.title characterizer
.include /home/shaheer/Desktop/FabRAM/FE/out/sram32x4.spi
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

      .tran 0.012144249999999999n 24.2885n 12.14425n
      .control
      set hcopydevtype = svg
      run
      meas tran tdiff_cell_rise TRIG v(clk) VAL=0.9 RISE=1 TARG v(Q0) VAL=0.9 RISE=1 
      meas tran tdiff_tran_rise TRIG v(Q0)  VAL=0.18000000000000002 RISE=1 TARG v(Q0) VAL=1.62 RISE=1 
      meas tran tdiff_cell_fall TRIG v(clk) VAL=0.9 RISE=2 TARG v(Q0) VAL=0.9 FALL=1 
      meas tran tdiff_tran_fall TRIG v(Q0)  VAL=1.62 FALL=1 TARG v(Q0) VAL=0.18000000000000002 FALL=1 

      echo "$&tdiff_cell_rise,$&tdiff_tran_rise $&tdiff_cell_fall,$&tdiff_tran_fall" > log/sim_0.42885_0.0379.text
      hardcopy log/sim_0.42885_0.0379.svg v(clk)+9.0 v(Q0)+7.2 v(x0.PCHG)+5.4 v(x0.WLEN)+3.6 v(x0.SAEN)+1.8 v(x0.WREN)
      exit
      .endc
      
Vpower VDD 0 1.8
Vgnd VSS 0 0
Vclk clk VSS DC 0V PULSE(0V 1.8V 0ns 0.5360625ns 0.5360625ns 2.5ns 6.072125ns)
Vaddr addr VSS DC 0V PULSE(0V 1.8V 0s 1ps 1ps 2.5ns 12.14425ns)
Vdin din VSS DC 0V PULSE(0V 1.8V 0s 1ps 1ps 2.5ns 12.14425ns)
Vwrite write VSS DC 0V PULSE(0V 1.8V 0s 1ps 1ps 12.14425ns 24.2885ns)
X0 VDD VSS clk addr addr addr addr addr din din din din Q0 Q1 Q2 Q3 write VDD sram32x4
C0 Q0 VSS 0.0379p
