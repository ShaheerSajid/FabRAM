magic
tech sky130A
magscale 1 2
timestamp 1702393006
<< nwell >>
rect 0 488 306 696
<< nmos >>
rect 94 201 124 285
rect 182 201 212 285
<< pmos >>
rect 94 550 124 634
rect 182 550 212 634
<< ndiff >>
rect 36 273 94 285
rect 36 213 48 273
rect 82 213 94 273
rect 36 201 94 213
rect 124 273 182 285
rect 124 213 136 273
rect 170 213 182 273
rect 124 201 182 213
rect 212 273 270 285
rect 212 213 224 273
rect 258 213 270 273
rect 212 201 270 213
<< pdiff >>
rect 36 622 94 634
rect 36 562 48 622
rect 82 562 94 622
rect 36 550 94 562
rect 124 622 182 634
rect 124 562 136 622
rect 170 562 182 622
rect 124 550 182 562
rect 212 622 270 634
rect 212 562 224 622
rect 258 562 270 622
rect 212 550 270 562
<< ndiffc >>
rect 48 213 82 273
rect 136 213 170 273
rect 224 213 258 273
<< pdiffc >>
rect 48 562 82 622
rect 136 562 170 622
rect 224 562 258 622
<< poly >>
rect 94 634 124 660
rect 182 634 212 660
rect 94 518 124 550
rect 44 502 124 518
rect 44 468 60 502
rect 94 468 124 502
rect 44 452 124 468
rect 94 285 124 452
rect 182 373 212 550
rect 182 357 262 373
rect 182 323 212 357
rect 246 323 262 357
rect 182 307 262 323
rect 182 285 212 307
rect 94 175 124 201
rect 182 175 212 201
<< polycont >>
rect 60 468 94 502
rect 212 323 246 357
<< locali >>
rect 48 622 82 638
rect 48 546 82 562
rect 136 622 170 638
rect 136 546 170 562
rect 224 622 258 638
rect 224 546 258 562
rect 44 468 60 502
rect 94 468 110 502
rect 48 323 60 357
rect 94 323 212 357
rect 246 323 262 357
rect 48 273 82 289
rect 48 197 82 213
rect 136 273 170 289
rect 136 197 170 213
rect 224 273 258 289
rect 224 197 258 213
<< viali >>
rect 48 562 82 622
rect 136 562 170 622
rect 224 562 258 622
rect 60 468 94 502
rect 60 323 94 357
rect 48 213 82 273
rect 136 213 170 273
rect 224 213 258 273
<< metal1 >>
rect 0 662 306 696
rect 48 634 82 662
rect 224 634 258 662
rect 42 622 88 634
rect 42 562 48 622
rect 82 562 88 622
rect 42 550 88 562
rect 130 622 176 634
rect 130 562 136 622
rect 170 562 176 622
rect 130 550 176 562
rect 218 622 264 634
rect 218 562 224 622
rect 258 562 264 622
rect 218 550 264 562
rect 48 502 106 508
rect 0 468 60 502
rect 94 468 106 502
rect 48 462 106 468
rect 136 444 170 550
rect 136 410 306 444
rect 48 357 106 363
rect 0 323 60 357
rect 94 323 106 357
rect 48 317 106 323
rect 136 285 170 410
rect 42 273 88 285
rect 42 213 48 273
rect 82 213 88 273
rect 42 201 88 213
rect 130 273 176 285
rect 130 213 136 273
rect 170 213 176 273
rect 130 201 176 213
rect 218 273 264 285
rect 218 213 224 273
rect 258 213 264 273
rect 218 201 264 213
rect 48 172 82 201
rect 224 172 258 201
rect 0 138 306 172
<< labels >>
rlabel metal1 0 662 34 696 0 VDD
rlabel metal1 0 468 34 502 0 A
rlabel metal1 0 323 34 357 0 B
rlabel metal1 0 138 34 172 0 VSS
rlabel metal1 272 410 306 444 0 Y
<< end >>
