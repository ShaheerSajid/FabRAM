magic
tech sky130A
magscale 1 2
timestamp 1703575910
<< nwell >>
rect 301 918 377 1126
rect 1013 1012 1184 1126
rect 1013 918 1043 1012
rect 1045 918 1168 1012
rect 1080 912 1298 918
rect 1655 917 1689 1126
rect 1080 521 1298 710
rect 1348 520 1437 521
rect 1348 312 1436 520
rect 1654 202 1688 521
rect 1772 234 1806 783
<< poly >>
rect 1130 932 1248 954
rect 1130 924 1172 932
rect 1156 898 1172 924
rect 1206 924 1248 932
rect 1206 898 1221 924
rect 1156 882 1221 898
rect 1173 876 1204 882
rect 65 312 95 349
rect -6 295 95 312
rect -6 261 11 295
rect 45 261 95 295
rect -6 245 95 261
rect 65 121 95 245
rect 283 209 313 349
rect 1782 231 1812 238
rect 2000 232 2030 238
rect 211 193 313 209
rect 211 159 227 193
rect 261 159 313 193
rect 1720 215 1812 231
rect 1720 181 1736 215
rect 1770 181 1812 215
rect 1720 165 1812 181
rect 1941 216 2030 232
rect 1941 182 1958 216
rect 1992 182 2030 216
rect 1941 166 2030 182
rect 211 143 313 159
rect 1782 152 1812 165
rect 2000 152 2030 166
rect 283 135 313 143
rect 1530 21 1560 34
rect 1468 5 1560 21
rect 1468 -29 1484 5
rect 1518 -29 1560 5
rect 1468 -45 1560 -29
rect 1530 -48 1560 -45
<< polycont >>
rect 1172 898 1206 932
rect 11 261 45 295
rect 227 159 261 193
rect 1736 181 1770 215
rect 1958 182 1992 216
rect 1484 -29 1518 5
<< locali >>
rect 1084 860 1118 976
rect 1156 898 1172 932
rect 1206 898 1390 932
rect 1084 854 1162 860
rect 1084 826 1152 854
rect 1356 806 1390 898
rect 323 753 425 787
rect 323 555 357 753
rect 107 521 357 555
rect 1574 547 1608 627
rect 107 463 141 521
rect 1374 513 1608 547
rect -6 261 11 295
rect 45 261 61 295
rect 107 193 141 371
rect 325 327 359 371
rect 325 293 450 327
rect 107 159 227 193
rect 261 159 277 193
rect 107 113 141 159
rect 325 113 359 293
rect 1374 182 1408 513
rect 1304 148 1408 182
rect 1699 181 1736 215
rect 1770 181 1786 215
rect 1824 130 1858 260
rect 1947 182 1958 216
rect 1992 182 2008 216
rect 2042 130 2076 260
rect 1266 5 1300 23
rect 1266 -29 1484 5
rect 1518 -29 1534 5
rect 1572 -70 1606 56
<< viali >>
rect 1356 772 1390 806
rect 11 261 45 295
rect 1665 181 1699 215
rect 1913 182 1947 216
<< metal1 >>
rect -1740 1092 -29 1126
rect 301 1092 377 1126
rect 1013 1092 1328 1126
rect 1354 1092 2124 1126
rect 1172 1064 1206 1092
rect 1736 1064 1770 1092
rect 1954 1064 1988 1092
rect 1026 992 1036 1044
rect 1089 992 1099 1044
rect 1290 992 1300 1044
rect 1353 992 1363 1044
rect 319 932 329 950
rect 273 898 329 932
rect 381 898 391 950
rect 273 880 301 898
rect 265 874 301 880
rect 1260 874 1294 980
rect -1740 840 -29 874
rect 273 870 301 874
rect 1013 678 1047 874
rect 1260 850 1326 874
rect 1232 840 1326 850
rect 1232 812 1294 840
rect 1344 806 1402 812
rect 1344 772 1356 806
rect 1390 802 1402 806
rect 1390 772 1636 802
rect 1344 766 1636 772
rect 1626 750 1636 766
rect 1688 750 1698 802
rect 1099 678 1109 730
rect -1740 568 -29 602
rect 301 568 377 602
rect 1013 568 1326 602
rect -1740 487 407 521
rect 1348 487 1730 521
rect 19 459 53 487
rect 237 459 271 487
rect 1484 458 1518 487
rect -1740 268 -218 302
rect -252 182 -218 268
rect -138 261 -128 313
rect -76 295 -66 313
rect -1 295 57 301
rect -76 261 11 295
rect 45 261 57 295
rect 1008 293 1042 326
rect 1008 281 1090 293
rect -1 255 57 261
rect 997 229 1007 281
rect 1059 229 1069 281
rect -252 148 406 182
rect 1648 175 1658 227
rect 1710 175 1720 227
rect 1762 172 1772 224
rect 1824 126 1858 264
rect 1894 175 1904 227
rect 1956 175 1966 227
rect 2042 126 2076 264
rect 2278 136 2576 145
rect 2278 84 2288 136
rect 2341 111 2576 136
rect 2341 84 2351 111
rect 19 -3 53 25
rect 237 -3 271 25
rect -1740 -37 444 -3
rect -138 -120 -128 -102
rect -1740 -154 -128 -120
rect -76 -154 -66 -102
rect 1348 -305 1382 -4
rect 1484 -305 1518 -274
rect 1736 -305 1770 -274
rect 1954 -305 1988 -274
rect 1348 -339 1988 -305
rect 2042 -589 2076 -274
rect 2042 -623 2576 -589
<< via1 >>
rect 1036 992 1089 1044
rect 1300 992 1353 1044
rect 329 898 381 950
rect 1636 750 1688 802
rect 1047 678 1099 730
rect -128 261 -76 313
rect 1007 229 1059 281
rect 1658 215 1710 227
rect 1658 181 1665 215
rect 1665 181 1699 215
rect 1699 181 1710 215
rect 1658 175 1710 181
rect 1772 172 1824 224
rect 1904 216 1956 227
rect 1904 182 1913 216
rect 1913 182 1947 216
rect 1947 182 1956 216
rect 1904 175 1956 182
rect 2288 84 2341 136
rect -128 -154 -76 -102
<< metal2 >>
rect 1025 1404 1077 1510
rect 918 1370 1077 1404
rect 918 1209 952 1370
rect 1894 1286 1946 1510
rect 55 1175 952 1209
rect 1055 1252 1946 1286
rect 1055 1178 1090 1252
rect 2484 1212 2536 1510
rect 1319 1178 2536 1212
rect -128 313 -76 323
rect -128 -102 -76 261
rect 55 253 89 1175
rect 1055 1054 1089 1178
rect 1319 1054 1353 1178
rect 1036 1044 1089 1054
rect 1036 982 1089 992
rect 1300 1044 1353 1054
rect 1300 982 1353 992
rect 329 950 381 960
rect 329 889 381 898
rect 329 854 1904 889
rect 1636 802 1688 812
rect 1688 750 1806 783
rect 1636 740 1806 750
rect 1047 730 1099 740
rect 1099 678 1658 702
rect 1047 668 1658 678
rect 1007 281 1059 291
rect 55 229 1007 253
rect 55 219 1059 229
rect 1624 237 1658 668
rect 1624 227 1710 237
rect 1624 175 1658 227
rect 1624 165 1710 175
rect 1772 234 1806 740
rect 1870 237 1904 854
rect 1772 224 1824 234
rect 1772 162 1824 172
rect 1870 227 1956 237
rect 1870 175 1904 227
rect 1870 165 1956 175
rect 1772 118 1806 162
rect 2288 136 2341 146
rect 1772 84 2288 118
rect 2288 74 2341 84
rect -128 -164 -76 -154
use sky130_fd_pr__nfet_01v8_A6LSUL  m1
timestamp 1703058996
transform 1 0 80 0 1 67
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m2
timestamp 1703056510
transform 1 0 80 0 1 417
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_A6LSUL  m3
timestamp 1703058996
transform 1 0 298 0 1 67
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m4
timestamp 1703056510
transform 1 0 298 0 1 417
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m5
timestamp 1703056510
transform 1 0 1189 0 1 808
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_54MHNA  m6
timestamp 1703060231
transform 1 0 1797 0 1 664
box -109 -462 109 462
use sky130_fd_pr__nfet_01v8_JB3UY8  m7
timestamp 1703060231
transform 1 0 1797 0 1 -74
box -73 -226 73 226
use sky130_fd_pr__pfet_01v8_54MHNA  m8
timestamp 1703060231
transform 1 0 2015 0 1 664
box -109 -462 109 462
use sky130_fd_pr__nfet_01v8_JB3UY8  m9
timestamp 1703060231
transform 1 0 2015 0 1 -74
box -73 -226 73 226
use nand2_f  nand2_f_0 ~/Desktop/FabRAM/FE/sram130/nand2
timestamp 1702829829
transform 1 0 406 0 1 -175
box 0 138 306 696
use nand2_f  nand2_f_1
timestamp 1702829829
transform 1 0 1042 0 1 -175
box 0 138 306 696
use nand2_f  nand2_f_2
timestamp 1702829829
transform 1 0 377 0 1 430
box 0 138 306 696
use not_f  not_f_0 ~/Desktop/FabRAM/FE/sram130/not
timestamp 1702826916
transform 1 0 712 0 1 -175
box 0 138 330 696
use not_f  not_f_1
timestamp 1702826916
transform 1 0 -29 0 1 430
box 0 138 330 696
use not_f  not_f_2
timestamp 1702826916
transform 1 0 683 0 1 430
box 0 138 330 696
use not_f  not_f_3
timestamp 1702826916
transform 1 0 1326 0 1 430
box 0 138 330 696
use sky130_fd_pr__nfet_01v8_L8ATA9  sky130_fd_pr__nfet_01v8_L8ATA9_0
timestamp 1703055308
transform 1 0 1545 0 1 -174
box -73 -126 73 126
use sky130_fd_pr__pfet_01v8_4Y88KP  sky130_fd_pr__pfet_01v8_4Y88KP_0
timestamp 1703056510
transform -1 0 1145 0 1 1022
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  sky130_fd_pr__pfet_01v8_4Y88KP_1
timestamp 1703056510
transform 1 0 1233 0 1 1022
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_5YUHNA  sky130_fd_pr__pfet_01v8_5YUHNA_0
timestamp 1703055308
transform 1 0 1545 0 1 259
box -109 -262 109 262
<< end >>
