magic
tech sky130A
magscale 1 2
timestamp 1702830205
<< nwell >>
rect 709 2146 1345 2354
rect 0 1560 1345 1768
rect 0 950 1345 1158
rect 709 360 1345 568
<< nmos >>
rect 803 1859 833 1943
rect 891 1859 921 1943
rect 1221 1859 1251 1943
rect 206 1273 236 1357
rect 803 1273 833 1357
rect 891 1273 921 1357
rect 1221 1273 1251 1357
rect 206 663 236 747
rect 803 663 833 747
rect 891 663 921 747
rect 1221 663 1251 747
rect 803 73 833 157
rect 891 73 921 157
rect 1221 73 1251 157
<< pmos >>
rect 803 2208 833 2292
rect 891 2208 921 2292
rect 1221 2208 1251 2292
rect 206 1622 236 1706
rect 803 1622 833 1706
rect 891 1622 921 1706
rect 1221 1622 1251 1706
rect 206 1012 236 1096
rect 803 1012 833 1096
rect 891 1012 921 1096
rect 1221 1012 1251 1096
rect 803 422 833 506
rect 891 422 921 506
rect 1221 422 1251 506
<< ndiff >>
rect 745 1931 803 1943
rect 745 1871 757 1931
rect 791 1871 803 1931
rect 745 1859 803 1871
rect 833 1931 891 1943
rect 833 1871 845 1931
rect 879 1871 891 1931
rect 833 1859 891 1871
rect 921 1931 979 1943
rect 921 1871 933 1931
rect 967 1871 979 1931
rect 921 1859 979 1871
rect 1163 1931 1221 1943
rect 1163 1871 1175 1931
rect 1209 1871 1221 1931
rect 1163 1859 1221 1871
rect 1251 1931 1309 1943
rect 1251 1871 1263 1931
rect 1297 1871 1309 1931
rect 1251 1859 1309 1871
rect 148 1345 206 1357
rect 148 1285 160 1345
rect 194 1285 206 1345
rect 148 1273 206 1285
rect 236 1345 294 1357
rect 236 1285 248 1345
rect 282 1285 294 1345
rect 236 1273 294 1285
rect 745 1345 803 1357
rect 745 1285 757 1345
rect 791 1285 803 1345
rect 745 1273 803 1285
rect 833 1345 891 1357
rect 833 1285 845 1345
rect 879 1285 891 1345
rect 833 1273 891 1285
rect 921 1345 979 1357
rect 921 1285 933 1345
rect 967 1285 979 1345
rect 921 1273 979 1285
rect 1163 1345 1221 1357
rect 1163 1285 1175 1345
rect 1209 1285 1221 1345
rect 1163 1273 1221 1285
rect 1251 1345 1309 1357
rect 1251 1285 1263 1345
rect 1297 1285 1309 1345
rect 1251 1273 1309 1285
rect 148 735 206 747
rect 148 675 160 735
rect 194 675 206 735
rect 148 663 206 675
rect 236 735 294 747
rect 236 675 248 735
rect 282 675 294 735
rect 236 663 294 675
rect 745 735 803 747
rect 745 675 757 735
rect 791 675 803 735
rect 745 663 803 675
rect 833 735 891 747
rect 833 675 845 735
rect 879 675 891 735
rect 833 663 891 675
rect 921 735 979 747
rect 921 675 933 735
rect 967 675 979 735
rect 921 663 979 675
rect 1163 735 1221 747
rect 1163 675 1175 735
rect 1209 675 1221 735
rect 1163 663 1221 675
rect 1251 735 1309 747
rect 1251 675 1263 735
rect 1297 675 1309 735
rect 1251 663 1309 675
rect 745 145 803 157
rect 745 85 757 145
rect 791 85 803 145
rect 745 73 803 85
rect 833 145 891 157
rect 833 85 845 145
rect 879 85 891 145
rect 833 73 891 85
rect 921 145 979 157
rect 921 85 933 145
rect 967 85 979 145
rect 921 73 979 85
rect 1163 145 1221 157
rect 1163 85 1175 145
rect 1209 85 1221 145
rect 1163 73 1221 85
rect 1251 145 1309 157
rect 1251 85 1263 145
rect 1297 85 1309 145
rect 1251 73 1309 85
<< pdiff >>
rect 745 2280 803 2292
rect 745 2220 757 2280
rect 791 2220 803 2280
rect 745 2208 803 2220
rect 833 2280 891 2292
rect 833 2220 845 2280
rect 879 2220 891 2280
rect 833 2208 891 2220
rect 921 2280 979 2292
rect 921 2220 933 2280
rect 967 2220 979 2280
rect 921 2208 979 2220
rect 1163 2280 1221 2292
rect 1163 2220 1175 2280
rect 1209 2220 1221 2280
rect 1163 2208 1221 2220
rect 1251 2280 1309 2292
rect 1251 2220 1263 2280
rect 1297 2220 1309 2280
rect 1251 2208 1309 2220
rect 148 1694 206 1706
rect 148 1634 160 1694
rect 194 1634 206 1694
rect 148 1622 206 1634
rect 236 1694 294 1706
rect 236 1634 248 1694
rect 282 1634 294 1694
rect 236 1622 294 1634
rect 745 1694 803 1706
rect 745 1634 757 1694
rect 791 1634 803 1694
rect 745 1622 803 1634
rect 833 1694 891 1706
rect 833 1634 845 1694
rect 879 1634 891 1694
rect 833 1622 891 1634
rect 921 1694 979 1706
rect 921 1634 933 1694
rect 967 1634 979 1694
rect 921 1622 979 1634
rect 1163 1694 1221 1706
rect 1163 1634 1175 1694
rect 1209 1634 1221 1694
rect 1163 1622 1221 1634
rect 1251 1694 1309 1706
rect 1251 1634 1263 1694
rect 1297 1634 1309 1694
rect 1251 1622 1309 1634
rect 148 1084 206 1096
rect 148 1024 160 1084
rect 194 1024 206 1084
rect 148 1012 206 1024
rect 236 1084 294 1096
rect 236 1024 248 1084
rect 282 1024 294 1084
rect 236 1012 294 1024
rect 745 1084 803 1096
rect 745 1024 757 1084
rect 791 1024 803 1084
rect 745 1012 803 1024
rect 833 1084 891 1096
rect 833 1024 845 1084
rect 879 1024 891 1084
rect 833 1012 891 1024
rect 921 1084 979 1096
rect 921 1024 933 1084
rect 967 1024 979 1084
rect 921 1012 979 1024
rect 1163 1084 1221 1096
rect 1163 1024 1175 1084
rect 1209 1024 1221 1084
rect 1163 1012 1221 1024
rect 1251 1084 1309 1096
rect 1251 1024 1263 1084
rect 1297 1024 1309 1084
rect 1251 1012 1309 1024
rect 745 494 803 506
rect 745 434 757 494
rect 791 434 803 494
rect 745 422 803 434
rect 833 494 891 506
rect 833 434 845 494
rect 879 434 891 494
rect 833 422 891 434
rect 921 494 979 506
rect 921 434 933 494
rect 967 434 979 494
rect 921 422 979 434
rect 1163 494 1221 506
rect 1163 434 1175 494
rect 1209 434 1221 494
rect 1163 422 1221 434
rect 1251 494 1309 506
rect 1251 434 1263 494
rect 1297 434 1309 494
rect 1251 422 1309 434
<< ndiffc >>
rect 757 1871 791 1931
rect 845 1871 879 1931
rect 933 1871 967 1931
rect 1175 1871 1209 1931
rect 1263 1871 1297 1931
rect 160 1285 194 1345
rect 248 1285 282 1345
rect 757 1285 791 1345
rect 845 1285 879 1345
rect 933 1285 967 1345
rect 1175 1285 1209 1345
rect 1263 1285 1297 1345
rect 160 675 194 735
rect 248 675 282 735
rect 757 675 791 735
rect 845 675 879 735
rect 933 675 967 735
rect 1175 675 1209 735
rect 1263 675 1297 735
rect 757 85 791 145
rect 845 85 879 145
rect 933 85 967 145
rect 1175 85 1209 145
rect 1263 85 1297 145
<< pdiffc >>
rect 757 2220 791 2280
rect 845 2220 879 2280
rect 933 2220 967 2280
rect 1175 2220 1209 2280
rect 1263 2220 1297 2280
rect 160 1634 194 1694
rect 248 1634 282 1694
rect 757 1634 791 1694
rect 845 1634 879 1694
rect 933 1634 967 1694
rect 1175 1634 1209 1694
rect 1263 1634 1297 1694
rect 160 1024 194 1084
rect 248 1024 282 1084
rect 757 1024 791 1084
rect 845 1024 879 1084
rect 933 1024 967 1084
rect 1175 1024 1209 1084
rect 1263 1024 1297 1084
rect 757 434 791 494
rect 845 434 879 494
rect 933 434 967 494
rect 1175 434 1209 494
rect 1263 434 1297 494
<< psubdiff >>
rect 1051 1931 1109 1955
rect 1051 1871 1063 1931
rect 1097 1871 1109 1931
rect 1051 1847 1109 1871
rect 36 1345 94 1369
rect 36 1285 48 1345
rect 82 1285 94 1345
rect 36 1261 94 1285
rect 1051 1345 1109 1369
rect 1051 1285 1063 1345
rect 1097 1285 1109 1345
rect 1051 1261 1109 1285
rect 36 735 94 759
rect 36 675 48 735
rect 82 675 94 735
rect 36 651 94 675
rect 1051 735 1109 759
rect 1051 675 1063 735
rect 1097 675 1109 735
rect 1051 651 1109 675
rect 1051 145 1109 169
rect 1051 85 1063 145
rect 1097 85 1109 145
rect 1051 61 1109 85
<< nsubdiff >>
rect 1051 2280 1109 2304
rect 1051 2220 1063 2280
rect 1097 2220 1109 2280
rect 1051 2196 1109 2220
rect 36 1694 94 1718
rect 36 1634 48 1694
rect 82 1634 94 1694
rect 36 1610 94 1634
rect 1051 1694 1109 1718
rect 1051 1634 1063 1694
rect 1097 1634 1109 1694
rect 1051 1610 1109 1634
rect 36 1084 94 1108
rect 36 1024 48 1084
rect 82 1024 94 1084
rect 36 1000 94 1024
rect 1051 1084 1109 1108
rect 1051 1024 1063 1084
rect 1097 1024 1109 1084
rect 1051 1000 1109 1024
rect 1051 494 1109 518
rect 1051 434 1063 494
rect 1097 434 1109 494
rect 1051 410 1109 434
<< psubdiffcont >>
rect 1063 1871 1097 1931
rect 48 1285 82 1345
rect 1063 1285 1097 1345
rect 48 675 82 735
rect 1063 675 1097 735
rect 1063 85 1097 145
<< nsubdiffcont >>
rect 1063 2220 1097 2280
rect 48 1634 82 1694
rect 1063 1634 1097 1694
rect 48 1024 82 1084
rect 1063 1024 1097 1084
rect 1063 434 1097 494
<< poly >>
rect 803 2292 833 2318
rect 891 2292 921 2318
rect 1221 2292 1251 2318
rect 803 2176 833 2208
rect 753 2160 833 2176
rect 753 2126 769 2160
rect 803 2126 833 2160
rect 753 2110 833 2126
rect 803 1943 833 2110
rect 891 2031 921 2208
rect 1221 2118 1251 2208
rect 1160 2102 1251 2118
rect 1160 2068 1176 2102
rect 1210 2068 1251 2102
rect 1160 2052 1251 2068
rect 891 2015 971 2031
rect 891 1981 921 2015
rect 955 1981 971 2015
rect 891 1965 971 1981
rect 891 1943 921 1965
rect 1221 1943 1251 2052
rect 803 1833 833 1859
rect 891 1833 921 1859
rect 1221 1833 1251 1859
rect 206 1706 236 1732
rect 803 1706 833 1732
rect 891 1706 921 1732
rect 1221 1706 1251 1732
rect 206 1532 236 1622
rect 803 1590 833 1622
rect 145 1516 236 1532
rect 753 1574 833 1590
rect 753 1540 769 1574
rect 803 1540 833 1574
rect 753 1524 833 1540
rect 145 1482 161 1516
rect 195 1482 236 1516
rect 145 1466 236 1482
rect 206 1357 236 1466
rect 803 1357 833 1524
rect 891 1445 921 1622
rect 1221 1532 1251 1622
rect 1160 1516 1251 1532
rect 1160 1482 1176 1516
rect 1210 1482 1251 1516
rect 1160 1466 1251 1482
rect 891 1429 971 1445
rect 891 1395 921 1429
rect 955 1395 971 1429
rect 891 1379 971 1395
rect 891 1357 921 1379
rect 1221 1357 1251 1466
rect 206 1247 236 1273
rect 803 1247 833 1273
rect 891 1247 921 1273
rect 1221 1247 1251 1273
rect 206 1096 236 1122
rect 803 1096 833 1122
rect 891 1096 921 1122
rect 1221 1096 1251 1122
rect 206 922 236 1012
rect 803 980 833 1012
rect 145 906 236 922
rect 753 964 833 980
rect 753 930 769 964
rect 803 930 833 964
rect 753 914 833 930
rect 145 872 161 906
rect 195 872 236 906
rect 145 856 236 872
rect 206 747 236 856
rect 803 747 833 914
rect 891 835 921 1012
rect 1221 922 1251 1012
rect 1160 906 1251 922
rect 1160 872 1176 906
rect 1210 872 1251 906
rect 1160 856 1251 872
rect 891 819 971 835
rect 891 785 921 819
rect 955 785 971 819
rect 891 769 971 785
rect 891 747 921 769
rect 1221 747 1251 856
rect 206 637 236 663
rect 803 637 833 663
rect 891 637 921 663
rect 1221 637 1251 663
rect 803 506 833 532
rect 891 506 921 532
rect 1221 506 1251 532
rect 803 390 833 422
rect 753 374 833 390
rect 753 340 769 374
rect 803 340 833 374
rect 753 324 833 340
rect 803 157 833 324
rect 891 245 921 422
rect 1221 332 1251 422
rect 1160 316 1251 332
rect 1160 282 1176 316
rect 1210 282 1251 316
rect 1160 266 1251 282
rect 891 229 971 245
rect 891 195 921 229
rect 955 195 971 229
rect 891 179 971 195
rect 891 157 921 179
rect 1221 157 1251 266
rect 803 47 833 73
rect 891 47 921 73
rect 1221 47 1251 73
<< polycont >>
rect 769 2126 803 2160
rect 1176 2068 1210 2102
rect 921 1981 955 2015
rect 769 1540 803 1574
rect 161 1482 195 1516
rect 1176 1482 1210 1516
rect 921 1395 955 1429
rect 769 930 803 964
rect 161 872 195 906
rect 1176 872 1210 906
rect 921 785 955 819
rect 769 340 803 374
rect 1176 282 1210 316
rect 921 195 955 229
<< locali >>
rect 757 2280 791 2296
rect 757 2204 791 2220
rect 845 2280 879 2296
rect 845 2204 879 2220
rect 933 2280 967 2296
rect 933 2204 967 2220
rect 1051 2280 1209 2296
rect 1051 2220 1063 2280
rect 1097 2220 1175 2280
rect 1051 2204 1209 2220
rect 1263 2280 1297 2296
rect 753 2126 769 2160
rect 803 2126 819 2160
rect 1263 2102 1297 2220
rect 1160 2068 1176 2102
rect 1210 2068 1226 2102
rect 757 1981 769 2015
rect 803 1981 921 2015
rect 955 1981 971 2015
rect 757 1931 791 1947
rect 757 1855 791 1871
rect 845 1931 879 1947
rect 845 1855 879 1871
rect 933 1931 967 1947
rect 933 1855 967 1871
rect 1063 1931 1209 1947
rect 1097 1871 1175 1931
rect 1063 1855 1209 1871
rect 1263 1931 1297 2068
rect 1263 1855 1297 1871
rect 36 1694 194 1710
rect 36 1634 48 1694
rect 82 1634 160 1694
rect 36 1618 194 1634
rect 248 1694 282 1710
rect 248 1516 282 1634
rect 757 1694 791 1710
rect 757 1618 791 1634
rect 845 1694 879 1710
rect 845 1618 879 1634
rect 933 1694 967 1710
rect 933 1618 967 1634
rect 1051 1694 1209 1710
rect 1051 1634 1063 1694
rect 1097 1634 1175 1694
rect 1051 1618 1209 1634
rect 1263 1694 1297 1710
rect 753 1540 769 1574
rect 803 1540 819 1574
rect 1263 1516 1297 1634
rect 145 1482 161 1516
rect 195 1482 211 1516
rect 1160 1482 1176 1516
rect 1210 1482 1226 1516
rect 48 1345 194 1361
rect 82 1285 160 1345
rect 48 1269 194 1285
rect 248 1345 282 1482
rect 757 1395 769 1429
rect 803 1395 921 1429
rect 955 1395 971 1429
rect 248 1269 282 1285
rect 757 1345 791 1361
rect 757 1269 791 1285
rect 845 1345 879 1361
rect 845 1269 879 1285
rect 933 1345 967 1361
rect 933 1269 967 1285
rect 1063 1345 1209 1361
rect 1097 1285 1175 1345
rect 1063 1269 1209 1285
rect 1263 1345 1297 1482
rect 1263 1269 1297 1285
rect 36 1084 194 1100
rect 36 1024 48 1084
rect 82 1024 160 1084
rect 36 1008 194 1024
rect 248 1084 282 1100
rect 248 906 282 1024
rect 757 1084 791 1100
rect 757 1008 791 1024
rect 845 1084 879 1100
rect 845 1008 879 1024
rect 933 1084 967 1100
rect 933 1008 967 1024
rect 1051 1084 1209 1100
rect 1051 1024 1063 1084
rect 1097 1024 1175 1084
rect 1051 1008 1209 1024
rect 1263 1084 1297 1100
rect 753 930 769 964
rect 803 930 819 964
rect 1263 906 1297 1024
rect 145 872 161 906
rect 195 872 211 906
rect 1160 872 1176 906
rect 1210 872 1226 906
rect 48 735 194 751
rect 82 675 160 735
rect 48 659 194 675
rect 248 735 282 872
rect 757 785 769 819
rect 803 785 921 819
rect 955 785 971 819
rect 248 659 282 675
rect 757 735 791 751
rect 757 659 791 675
rect 845 735 879 751
rect 845 659 879 675
rect 933 735 967 751
rect 933 659 967 675
rect 1063 735 1209 751
rect 1097 675 1175 735
rect 1063 659 1209 675
rect 1263 735 1297 872
rect 1263 659 1297 675
rect 757 494 791 510
rect 757 418 791 434
rect 845 494 879 510
rect 845 418 879 434
rect 933 494 967 510
rect 933 418 967 434
rect 1051 494 1209 510
rect 1051 434 1063 494
rect 1097 434 1175 494
rect 1051 418 1209 434
rect 1263 494 1297 510
rect 753 340 769 374
rect 803 340 819 374
rect 1263 316 1297 434
rect 1160 282 1176 316
rect 1210 282 1226 316
rect 757 195 769 229
rect 803 195 921 229
rect 955 195 971 229
rect 757 145 791 161
rect 757 69 791 85
rect 845 145 879 161
rect 845 69 879 85
rect 933 145 967 161
rect 933 69 967 85
rect 1063 145 1209 161
rect 1097 85 1175 145
rect 1063 69 1209 85
rect 1263 145 1297 282
rect 1263 69 1297 85
<< viali >>
rect 757 2220 791 2280
rect 845 2220 879 2280
rect 933 2220 967 2280
rect 1175 2220 1209 2280
rect 1263 2220 1297 2280
rect 769 2126 803 2160
rect 1176 2068 1210 2102
rect 1263 2068 1297 2102
rect 769 1981 803 2015
rect 757 1871 791 1931
rect 845 1871 879 1931
rect 933 1871 967 1931
rect 1175 1871 1209 1931
rect 1263 1871 1297 1931
rect 160 1634 194 1694
rect 248 1634 282 1694
rect 757 1634 791 1694
rect 845 1634 879 1694
rect 933 1634 967 1694
rect 1175 1634 1209 1694
rect 1263 1634 1297 1694
rect 769 1540 803 1574
rect 161 1482 195 1516
rect 248 1482 282 1516
rect 1176 1482 1210 1516
rect 1263 1482 1297 1516
rect 160 1285 194 1345
rect 769 1395 803 1429
rect 248 1285 282 1345
rect 757 1285 791 1345
rect 845 1285 879 1345
rect 933 1285 967 1345
rect 1175 1285 1209 1345
rect 1263 1285 1297 1345
rect 160 1024 194 1084
rect 248 1024 282 1084
rect 757 1024 791 1084
rect 845 1024 879 1084
rect 933 1024 967 1084
rect 1175 1024 1209 1084
rect 1263 1024 1297 1084
rect 769 930 803 964
rect 161 872 195 906
rect 248 872 282 906
rect 1176 872 1210 906
rect 1263 872 1297 906
rect 160 675 194 735
rect 769 785 803 819
rect 248 675 282 735
rect 757 675 791 735
rect 845 675 879 735
rect 933 675 967 735
rect 1175 675 1209 735
rect 1263 675 1297 735
rect 757 434 791 494
rect 845 434 879 494
rect 933 434 967 494
rect 1175 434 1209 494
rect 1263 434 1297 494
rect 769 340 803 374
rect 1176 282 1210 316
rect 1263 282 1297 316
rect 769 195 803 229
rect 757 85 791 145
rect 845 85 879 145
rect 933 85 967 145
rect 1175 85 1209 145
rect 1263 85 1297 145
<< metal1 >>
rect 637 2302 647 2354
rect 699 2320 1345 2354
rect 699 2302 709 2320
rect 757 2292 791 2320
rect 933 2292 967 2320
rect 1175 2292 1209 2320
rect 751 2280 797 2292
rect 751 2220 757 2280
rect 791 2220 797 2280
rect 751 2208 797 2220
rect 839 2280 885 2292
rect 839 2220 845 2280
rect 879 2220 885 2280
rect 839 2208 885 2220
rect 927 2280 973 2292
rect 927 2220 933 2280
rect 967 2220 973 2280
rect 927 2208 973 2220
rect 1169 2280 1215 2292
rect 1169 2220 1175 2280
rect 1209 2220 1215 2280
rect 1169 2208 1215 2220
rect 1257 2280 1303 2292
rect 1257 2220 1263 2280
rect 1297 2220 1303 2280
rect 1257 2208 1303 2220
rect 477 2126 487 2178
rect 539 2160 549 2178
rect 757 2160 815 2166
rect 539 2126 769 2160
rect 803 2126 815 2160
rect 757 2120 815 2126
rect 845 2102 879 2208
rect 1299 2108 1309 2111
rect 1164 2102 1222 2108
rect 845 2068 1176 2102
rect 1210 2068 1222 2102
rect 397 1981 407 2033
rect 459 2015 469 2033
rect 757 2015 815 2021
rect 459 1981 769 2015
rect 803 1981 815 2015
rect 757 1975 815 1981
rect 933 1943 967 2068
rect 1164 2062 1222 2068
rect 1251 2102 1309 2108
rect 1251 2068 1263 2102
rect 1297 2068 1309 2102
rect 1251 2062 1309 2068
rect 1299 2059 1309 2062
rect 1361 2059 1371 2111
rect 751 1931 797 1943
rect 751 1871 757 1931
rect 791 1871 797 1931
rect 751 1859 797 1871
rect 839 1931 885 1943
rect 839 1871 845 1931
rect 879 1871 885 1931
rect 839 1859 885 1871
rect 927 1931 973 1943
rect 927 1871 933 1931
rect 967 1871 973 1931
rect 927 1859 973 1871
rect 1169 1931 1215 1943
rect 1169 1871 1175 1931
rect 1209 1871 1215 1931
rect 1169 1859 1215 1871
rect 1257 1931 1303 1943
rect 1257 1871 1263 1931
rect 1297 1871 1303 1931
rect 1257 1859 1303 1871
rect 557 1796 567 1848
rect 619 1830 629 1848
rect 757 1830 791 1859
rect 1175 1830 1209 1859
rect 619 1796 1345 1830
rect 0 1734 647 1768
rect 160 1706 194 1734
rect 637 1716 647 1734
rect 699 1734 1345 1768
rect 699 1716 709 1734
rect 757 1706 791 1734
rect 933 1706 967 1734
rect 1175 1706 1209 1734
rect 154 1694 200 1706
rect 154 1634 160 1694
rect 194 1634 200 1694
rect 154 1622 200 1634
rect 242 1694 288 1706
rect 242 1634 248 1694
rect 282 1634 288 1694
rect 242 1622 288 1634
rect 751 1694 797 1706
rect 751 1634 757 1694
rect 791 1634 797 1694
rect 751 1622 797 1634
rect 839 1694 885 1706
rect 839 1634 845 1694
rect 879 1634 885 1694
rect 839 1622 885 1634
rect 927 1694 973 1706
rect 927 1634 933 1694
rect 967 1634 973 1694
rect 927 1622 973 1634
rect 1169 1694 1215 1706
rect 1169 1634 1175 1694
rect 1209 1634 1215 1694
rect 1169 1622 1215 1634
rect 1257 1694 1303 1706
rect 1257 1634 1263 1694
rect 1297 1634 1303 1694
rect 1257 1622 1303 1634
rect 477 1540 487 1592
rect 539 1574 549 1592
rect 757 1574 815 1580
rect 539 1540 769 1574
rect 803 1540 815 1574
rect 149 1516 207 1522
rect 0 1482 161 1516
rect 195 1482 207 1516
rect 149 1476 207 1482
rect 236 1516 294 1522
rect 477 1516 505 1540
rect 757 1534 815 1540
rect 236 1482 248 1516
rect 282 1482 505 1516
rect 845 1516 879 1622
rect 1299 1522 1309 1525
rect 1164 1516 1222 1522
rect 845 1482 1176 1516
rect 1210 1482 1222 1516
rect 236 1476 294 1482
rect 161 1439 195 1476
rect 477 1439 487 1448
rect 161 1405 487 1439
rect 477 1396 487 1405
rect 539 1396 549 1448
rect 757 1429 815 1435
rect 647 1395 769 1429
rect 803 1395 815 1429
rect 154 1345 200 1357
rect 154 1285 160 1345
rect 194 1285 200 1345
rect 154 1273 200 1285
rect 242 1345 288 1357
rect 242 1285 248 1345
rect 282 1285 288 1345
rect 317 1310 327 1362
rect 379 1344 389 1362
rect 647 1344 681 1395
rect 757 1389 815 1395
rect 933 1357 967 1482
rect 1164 1476 1222 1482
rect 1251 1516 1309 1522
rect 1251 1482 1263 1516
rect 1297 1482 1309 1516
rect 1251 1476 1309 1482
rect 1299 1473 1309 1476
rect 1361 1473 1371 1525
rect 379 1310 681 1344
rect 751 1345 797 1357
rect 242 1273 288 1285
rect 751 1285 757 1345
rect 791 1285 797 1345
rect 751 1273 797 1285
rect 839 1345 885 1357
rect 839 1285 845 1345
rect 879 1285 885 1345
rect 839 1273 885 1285
rect 927 1345 973 1357
rect 927 1285 933 1345
rect 967 1285 973 1345
rect 927 1273 973 1285
rect 1169 1345 1215 1357
rect 1169 1285 1175 1345
rect 1209 1285 1215 1345
rect 1169 1273 1215 1285
rect 1257 1345 1303 1357
rect 1257 1285 1263 1345
rect 1297 1285 1303 1345
rect 1257 1273 1303 1285
rect 160 1244 194 1273
rect 557 1244 567 1272
rect 0 1220 567 1244
rect 619 1244 629 1272
rect 757 1244 791 1273
rect 1175 1244 1209 1273
rect 619 1220 1345 1244
rect 0 1210 1345 1220
rect 327 1209 455 1210
rect 0 1124 647 1158
rect 160 1096 194 1124
rect 637 1106 647 1124
rect 699 1124 1345 1158
rect 699 1106 709 1124
rect 757 1096 791 1124
rect 933 1096 967 1124
rect 1175 1096 1209 1124
rect 154 1084 200 1096
rect 154 1024 160 1084
rect 194 1024 200 1084
rect 154 1012 200 1024
rect 242 1084 288 1096
rect 242 1024 248 1084
rect 282 1024 288 1084
rect 242 1012 288 1024
rect 751 1084 797 1096
rect 751 1024 757 1084
rect 791 1024 797 1084
rect 751 1012 797 1024
rect 839 1084 885 1096
rect 839 1024 845 1084
rect 879 1024 885 1084
rect 839 1012 885 1024
rect 927 1084 973 1096
rect 927 1024 933 1084
rect 967 1024 973 1084
rect 927 1012 973 1024
rect 1169 1084 1215 1096
rect 1169 1024 1175 1084
rect 1209 1024 1215 1084
rect 1169 1012 1215 1024
rect 1257 1084 1303 1096
rect 1257 1024 1263 1084
rect 1297 1024 1303 1084
rect 1257 1012 1303 1024
rect 477 930 487 982
rect 539 964 549 982
rect 757 964 815 970
rect 539 930 769 964
rect 803 930 815 964
rect 757 924 815 930
rect 149 906 207 912
rect 0 872 161 906
rect 195 872 207 906
rect 149 866 207 872
rect 236 906 294 912
rect 845 906 879 1012
rect 1299 912 1309 915
rect 1164 906 1222 912
rect 236 872 248 906
rect 282 872 431 906
rect 845 872 1176 906
rect 1210 872 1222 906
rect 236 866 294 872
rect 161 811 195 866
rect 397 837 431 872
rect 161 777 351 811
rect 397 785 407 837
rect 459 819 469 837
rect 757 819 815 825
rect 459 785 769 819
rect 803 785 815 819
rect 757 779 815 785
rect 154 735 200 747
rect 154 675 160 735
rect 194 675 200 735
rect 154 663 200 675
rect 242 735 288 747
rect 242 675 248 735
rect 282 675 288 735
rect 317 734 351 777
rect 933 747 967 872
rect 1164 866 1222 872
rect 1251 906 1309 912
rect 1251 872 1263 906
rect 1297 872 1309 906
rect 1251 866 1309 872
rect 1299 863 1309 866
rect 1361 863 1371 915
rect 751 735 797 747
rect 317 682 327 734
rect 379 682 389 734
rect 242 663 288 675
rect 751 675 757 735
rect 791 675 797 735
rect 751 663 797 675
rect 839 735 885 747
rect 839 675 845 735
rect 879 675 885 735
rect 839 663 885 675
rect 927 735 973 747
rect 927 675 933 735
rect 967 675 973 735
rect 927 663 973 675
rect 1169 735 1215 747
rect 1169 675 1175 735
rect 1209 675 1215 735
rect 1169 663 1215 675
rect 1257 735 1303 747
rect 1257 675 1263 735
rect 1297 675 1303 735
rect 1257 663 1303 675
rect 160 634 194 663
rect 557 634 567 662
rect 0 610 567 634
rect 619 634 629 662
rect 757 634 791 663
rect 1175 634 1209 663
rect 619 610 1345 634
rect 0 600 1345 610
rect 637 516 647 568
rect 699 534 1345 568
rect 699 516 709 534
rect 757 506 791 534
rect 933 506 967 534
rect 1175 506 1209 534
rect 751 494 797 506
rect 751 434 757 494
rect 791 434 797 494
rect 751 422 797 434
rect 839 494 885 506
rect 839 434 845 494
rect 879 434 885 494
rect 839 422 885 434
rect 927 494 973 506
rect 927 434 933 494
rect 967 434 973 494
rect 927 422 973 434
rect 1169 494 1215 506
rect 1169 434 1175 494
rect 1209 434 1215 494
rect 1169 422 1215 434
rect 1257 494 1303 506
rect 1257 434 1263 494
rect 1297 434 1303 494
rect 1257 422 1303 434
rect 477 340 487 392
rect 539 374 549 392
rect 757 374 815 380
rect 539 340 769 374
rect 803 340 815 374
rect 757 334 815 340
rect 845 316 879 422
rect 1299 322 1309 325
rect 1164 316 1222 322
rect 845 282 1176 316
rect 1210 282 1222 316
rect 316 195 326 247
rect 378 229 388 247
rect 757 229 815 235
rect 378 195 769 229
rect 803 195 815 229
rect 757 189 815 195
rect 933 157 967 282
rect 1164 276 1222 282
rect 1251 316 1309 322
rect 1251 282 1263 316
rect 1297 282 1309 316
rect 1251 276 1309 282
rect 1299 273 1309 276
rect 1361 273 1371 325
rect 751 145 797 157
rect 751 85 757 145
rect 791 85 797 145
rect 751 73 797 85
rect 839 145 885 157
rect 839 85 845 145
rect 879 85 885 145
rect 839 73 885 85
rect 927 145 973 157
rect 927 85 933 145
rect 967 85 973 145
rect 927 73 973 85
rect 1169 145 1215 157
rect 1169 85 1175 145
rect 1209 85 1215 145
rect 1169 73 1215 85
rect 1257 145 1303 157
rect 1257 85 1263 145
rect 1297 85 1303 145
rect 1257 73 1303 85
rect 557 10 567 62
rect 619 44 629 62
rect 757 44 791 73
rect 1175 44 1209 73
rect 619 10 1345 44
<< via1 >>
rect 647 2302 699 2354
rect 487 2126 539 2178
rect 407 1981 459 2033
rect 1309 2059 1361 2111
rect 567 1796 619 1848
rect 647 1716 699 1768
rect 487 1540 539 1592
rect 487 1396 539 1448
rect 327 1310 379 1362
rect 1309 1473 1361 1525
rect 567 1220 619 1272
rect 647 1106 699 1158
rect 487 930 539 982
rect 407 785 459 837
rect 1309 863 1361 915
rect 327 682 379 734
rect 567 610 619 662
rect 647 516 699 568
rect 487 340 539 392
rect 326 195 378 247
rect 1309 273 1361 325
rect 567 10 619 62
<< metal2 >>
rect 487 2178 539 2188
rect 407 2033 459 2043
rect 327 1362 379 1372
rect 327 734 379 1310
rect 407 837 459 1981
rect 487 1592 539 2126
rect 487 1534 539 1540
rect 567 1848 619 2422
rect 407 777 459 785
rect 487 1448 539 1456
rect 487 982 539 1396
rect 327 257 379 682
rect 487 392 539 930
rect 487 331 539 340
rect 567 1272 619 1796
rect 567 662 619 1220
rect 326 247 379 257
rect 378 195 379 247
rect 326 185 379 195
rect 567 62 619 610
rect 567 0 619 10
rect 647 2354 699 2422
rect 647 1768 699 2302
rect 1307 2113 1363 2123
rect 1307 2047 1363 2057
rect 647 1158 699 1716
rect 1307 1527 1363 1537
rect 1307 1461 1363 1471
rect 647 568 699 1106
rect 1307 917 1363 927
rect 1307 851 1363 861
rect 647 0 699 516
rect 1307 327 1363 337
rect 1307 261 1363 271
<< via2 >>
rect 1307 2111 1363 2113
rect 1307 2059 1309 2111
rect 1309 2059 1361 2111
rect 1361 2059 1363 2111
rect 1307 2057 1363 2059
rect 1307 1525 1363 1527
rect 1307 1473 1309 1525
rect 1309 1473 1361 1525
rect 1361 1473 1363 1525
rect 1307 1471 1363 1473
rect 1307 915 1363 917
rect 1307 863 1309 915
rect 1309 863 1361 915
rect 1361 863 1363 915
rect 1307 861 1363 863
rect 1307 325 1363 327
rect 1307 273 1309 325
rect 1309 273 1361 325
rect 1361 273 1363 325
rect 1307 271 1363 273
<< metal3 >>
rect 1297 2113 1462 2118
rect 1297 2057 1307 2113
rect 1363 2057 1462 2113
rect 1297 2052 1462 2057
rect 1297 1527 1462 1532
rect 1297 1471 1307 1527
rect 1363 1471 1462 1527
rect 1297 1466 1462 1471
rect 1297 917 1462 922
rect 1297 861 1307 917
rect 1363 861 1462 917
rect 1297 856 1462 861
rect 1297 327 1462 332
rect 1297 271 1307 327
rect 1363 271 1462 327
rect 1297 266 1462 271
<< labels >>
rlabel metal3 1396 2052 1462 2118 0 Y0
rlabel metal3 1396 1466 1462 1532 0 Y1
rlabel metal3 1396 856 1462 922 0 Y2
rlabel metal3 1396 266 1462 332 0 Y3
rlabel metal2 567 2370 619 2422 0 VSS
rlabel metal2 647 2370 699 2422 0 VDD
rlabel metal1 0 1482 34 1516 0 A1
rlabel metal1 0 872 34 906 0 A0
<< end >>
