magic
tech sky130A
magscale 1 2
timestamp 1703664600
<< metal1 >>
rect 985 4916 995 4938
rect 831 4882 995 4916
rect 1051 4882 1061 4938
rect 1079 4220 1089 4242
rect 831 4186 1089 4220
rect 1145 4186 1155 4242
rect 1163 3524 1173 3546
rect 831 3490 1173 3524
rect 1229 3490 1239 3546
rect 2179 3389 2213 5275
rect 2179 3355 2289 3389
rect 1257 2828 1267 2850
rect 831 2794 1267 2828
rect 1323 2794 1333 2850
rect 1341 2132 1351 2154
rect 831 2098 1351 2132
rect 1407 2098 1417 2154
rect 1437 1436 1447 1458
rect 831 1402 1447 1436
rect 1503 1402 1513 1458
rect 1544 740 1554 762
rect 831 706 1554 740
rect 1610 706 1620 762
rect 1642 44 1652 66
rect 831 10 1652 44
rect 1708 10 1718 66
<< via1 >>
rect 995 4882 1051 4938
rect 1089 4186 1145 4242
rect 1173 3490 1229 3546
rect 1267 2794 1323 2850
rect 1351 2098 1407 2154
rect 1447 1402 1503 1458
rect 1554 706 1610 762
rect 1652 10 1708 66
<< metal2 >>
rect 0 5167 53 5275
rect 995 5145 1051 5155
rect 995 4938 1051 5089
rect 995 4872 1051 4882
rect 1089 5019 1145 5029
rect 1089 4242 1145 4963
rect 1089 4152 1145 4186
rect 1173 4893 1229 4903
rect 1173 3546 1229 4837
rect 1173 3472 1229 3490
rect 1267 4767 1323 4777
rect 1267 2850 1323 4711
rect 1267 2783 1323 2794
rect 1351 4641 1407 4651
rect 1351 4575 1407 4585
rect 1351 2164 1406 4575
rect 1447 4515 1503 4525
rect 1351 2154 1407 2164
rect 1351 2088 1407 2098
rect 1447 1458 1503 4459
rect 1447 1389 1503 1402
rect 1554 4389 1610 4399
rect 1554 762 1610 4333
rect 1554 696 1610 706
rect 1652 4263 1708 4273
rect 1652 66 1708 4207
rect 1652 0 1708 10
<< via2 >>
rect 995 5089 1051 5145
rect 1089 4963 1145 5019
rect 1173 4837 1229 4893
rect 1267 4711 1323 4767
rect 1351 4585 1407 4641
rect 1447 4459 1503 4515
rect 1554 4333 1610 4389
rect 1652 4207 1708 4263
<< metal3 >>
rect 985 5145 2289 5150
rect 985 5089 995 5145
rect 1051 5089 2289 5145
rect 985 5084 2289 5089
rect 1079 5019 2289 5024
rect 1079 4963 1089 5019
rect 1145 4963 2289 5019
rect 1079 4958 2289 4963
rect 1163 4893 2289 4898
rect 1163 4837 1173 4893
rect 1229 4837 2289 4893
rect 1163 4832 2289 4837
rect 1257 4767 2289 4772
rect 1257 4711 1267 4767
rect 1323 4711 2289 4767
rect 1257 4706 2289 4711
rect 1341 4641 2289 4646
rect 1341 4585 1351 4641
rect 1407 4585 2289 4641
rect 1341 4580 2289 4585
rect 1437 4515 2289 4520
rect 1437 4459 1447 4515
rect 1503 4459 2289 4515
rect 1437 4454 2289 4459
rect 1544 4389 2289 4394
rect 1544 4333 1554 4389
rect 1610 4333 2289 4389
rect 1544 4328 2289 4333
rect 1642 4263 2289 4268
rect 1642 4207 1652 4263
rect 1708 4207 2289 4263
rect 1642 4202 2289 4207
<< labels >>
rlabel metal1 831 4882 865 4916 0 SEL0
rlabel metal1 831 4186 865 4220 0 SEL1
rlabel metal1 831 3490 865 3524 0 SEL2
rlabel metal1 831 2794 865 2828 0 SEL3
rlabel metal1 831 2098 865 2132 0 SEL4
rlabel metal1 831 1402 865 1436 0 SEL5
rlabel metal1 831 706 865 740 0 SEL6
rlabel metal1 831 10 865 44 0 SEL7
<< end >>
