magic
tech sky130A
magscale 1 2
timestamp 1703662019
<< metal1 >>
rect 985 2133 995 2155
rect 831 2099 995 2133
rect 1051 2099 1061 2155
rect 1079 1437 1089 1459
rect 831 1403 1089 1437
rect 1145 1403 1155 1459
rect 2179 1110 2213 2492
rect 2179 1076 2300 1110
rect 1163 741 1173 763
rect 831 707 1173 741
rect 1229 707 1239 763
rect 1257 45 1267 67
rect 831 11 1267 45
rect 1323 11 1333 67
<< via1 >>
rect 995 2099 1051 2155
rect 1089 1403 1145 1459
rect 1173 707 1229 763
rect 1267 11 1323 67
<< metal2 >>
rect 0 2384 53 2492
rect 995 2362 1051 2372
rect 995 2155 1051 2306
rect 995 2089 1051 2099
rect 1089 2236 1145 2246
rect 1089 1459 1145 2180
rect 1089 1369 1145 1403
rect 1173 2110 1229 2120
rect 1173 763 1229 2054
rect 1173 689 1229 707
rect 1267 1984 1323 1994
rect 1267 67 1323 1928
rect 1267 0 1323 11
<< via2 >>
rect 995 2306 1051 2362
rect 1089 2180 1145 2236
rect 1173 2054 1229 2110
rect 1267 1928 1323 1984
<< metal3 >>
rect 985 2362 2289 2367
rect 985 2306 995 2362
rect 1051 2306 2289 2362
rect 985 2301 2289 2306
rect 1079 2236 2289 2241
rect 1079 2180 1089 2236
rect 1145 2180 2289 2236
rect 1079 2175 2289 2180
rect 1163 2110 2289 2115
rect 1163 2054 1173 2110
rect 1229 2054 2289 2110
rect 1163 2049 2289 2054
rect 1257 1984 2289 1989
rect 1257 1928 1267 1984
rect 1323 1928 2289 1984
rect 1257 1923 2289 1928
<< labels >>
rlabel metal1 831 2099 865 2133 0 SEL0
rlabel metal1 831 1403 865 1437 0 SEL1
rlabel metal1 831 707 865 741 0 SEL2
rlabel metal1 831 11 865 45 0 SEL3
<< end >>
