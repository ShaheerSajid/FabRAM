magic
tech sky130A
magscale 1 2
timestamp 1702386302
<< nwell >>
rect 0 488 720 696
<< nmos >>
rect 93 200 123 320
rect 293 200 323 360
rect 381 200 411 360
rect 595 200 625 320
<< pmos >>
rect 293 550 323 634
rect 381 550 411 634
<< ndiff >>
rect 235 348 293 360
rect 35 308 93 320
rect 35 212 47 308
rect 81 212 93 308
rect 35 200 93 212
rect 123 308 181 320
rect 123 212 135 308
rect 169 212 181 308
rect 123 200 181 212
rect 235 212 247 348
rect 281 212 293 348
rect 235 200 293 212
rect 323 348 381 360
rect 323 212 335 348
rect 369 212 381 348
rect 323 200 381 212
rect 411 348 469 360
rect 411 212 423 348
rect 457 212 469 348
rect 411 200 469 212
rect 537 308 595 320
rect 537 212 549 308
rect 583 212 595 308
rect 537 200 595 212
rect 625 308 683 320
rect 625 212 637 308
rect 671 212 683 308
rect 625 200 683 212
<< pdiff >>
rect 235 622 293 634
rect 235 562 247 622
rect 281 562 293 622
rect 235 550 293 562
rect 323 622 381 634
rect 323 562 335 622
rect 369 562 381 622
rect 323 550 381 562
rect 411 622 469 634
rect 411 562 423 622
rect 457 562 469 622
rect 411 550 469 562
<< ndiffc >>
rect 47 212 81 308
rect 135 212 169 308
rect 247 212 281 348
rect 335 212 369 348
rect 423 212 457 348
rect 549 212 583 308
rect 637 212 671 308
<< pdiffc >>
rect 247 562 281 622
rect 335 562 369 622
rect 423 562 457 622
<< psubdiff >>
rect 310 122 392 146
rect 310 88 335 122
rect 369 88 392 122
rect 310 64 392 88
<< nsubdiff >>
rect 523 622 605 634
rect 523 562 547 622
rect 581 562 605 622
rect 523 550 605 562
<< psubdiffcont >>
rect 335 88 369 122
<< nsubdiffcont >>
rect 547 562 581 622
<< poly >>
rect 293 634 323 660
rect 381 634 411 660
rect 293 515 323 550
rect 257 503 323 515
rect 257 469 273 503
rect 307 469 323 503
rect 257 458 323 469
rect 27 435 123 451
rect 27 401 43 435
rect 77 401 123 435
rect 27 385 123 401
rect 93 320 123 385
rect 293 360 323 458
rect 381 447 411 550
rect 381 432 447 447
rect 381 398 397 432
rect 431 398 447 432
rect 381 381 447 398
rect 578 435 644 451
rect 578 401 594 435
rect 628 401 644 435
rect 578 385 644 401
rect 381 360 411 381
rect 595 320 625 385
rect 93 174 123 200
rect 293 174 323 200
rect 381 174 411 200
rect 595 174 625 200
<< polycont >>
rect 273 469 307 503
rect 43 401 77 435
rect 397 398 431 432
rect 594 401 628 435
<< locali >>
rect 247 622 281 638
rect 189 562 247 580
rect 189 546 281 562
rect 335 622 369 638
rect 335 546 369 562
rect 423 622 457 638
rect 27 401 34 435
rect 86 401 93 435
rect 189 432 223 546
rect 423 503 457 562
rect 547 622 581 646
rect 547 538 581 562
rect 257 469 273 503
rect 307 469 515 503
rect 135 398 397 432
rect 431 398 447 432
rect 47 308 81 324
rect 47 196 81 212
rect 135 308 169 398
rect 135 196 169 212
rect 247 348 281 398
rect 481 364 515 469
rect 578 401 585 435
rect 637 401 644 435
rect 247 196 281 212
rect 335 348 369 364
rect 335 196 369 212
rect 423 348 583 364
rect 457 330 583 348
rect 423 196 457 212
rect 549 308 583 330
rect 549 196 583 212
rect 637 308 671 324
rect 637 196 671 212
rect 310 122 392 146
rect 310 88 335 122
rect 369 88 392 122
rect 310 64 392 88
<< viali >>
rect 247 562 281 622
rect 335 562 369 622
rect 423 562 457 622
rect 34 435 86 453
rect 34 401 43 435
rect 43 401 77 435
rect 77 401 86 435
rect 547 562 581 622
rect 47 212 81 308
rect 135 212 169 308
rect 585 435 637 453
rect 585 401 594 435
rect 594 401 628 435
rect 628 401 637 435
rect 247 212 281 348
rect 335 212 369 348
rect 423 212 457 348
rect 549 212 583 308
rect 637 212 671 308
rect 335 88 369 122
<< metal1 >>
rect 0 662 720 696
rect 335 634 369 662
rect 547 634 581 662
rect 241 622 287 634
rect 241 562 247 622
rect 281 562 287 622
rect 241 550 287 562
rect 329 622 375 634
rect 329 562 335 622
rect 369 562 375 622
rect 329 550 375 562
rect 417 622 463 634
rect 417 562 423 622
rect 457 562 463 622
rect 417 550 463 562
rect 541 622 587 634
rect 541 562 547 622
rect 581 562 587 622
rect 541 550 587 562
rect 22 453 98 459
rect 22 444 34 453
rect 0 410 34 444
rect 22 401 34 410
rect 86 444 98 453
rect 573 453 649 459
rect 573 444 585 453
rect 86 410 585 444
rect 86 401 98 410
rect 22 395 98 401
rect 573 401 585 410
rect 637 444 649 453
rect 637 410 720 444
rect 637 401 649 410
rect 573 395 649 401
rect 241 348 287 360
rect 41 308 87 320
rect 41 258 47 308
rect 81 258 87 308
rect 129 308 175 320
rect 28 206 38 258
rect 90 206 100 258
rect 129 212 135 308
rect 169 212 175 308
rect 41 200 87 206
rect 129 200 175 212
rect 241 212 247 348
rect 281 212 287 348
rect 241 200 287 212
rect 329 348 375 360
rect 329 212 335 348
rect 369 212 375 348
rect 329 200 375 212
rect 417 348 463 360
rect 417 212 423 348
rect 457 212 463 348
rect 417 200 463 212
rect 543 308 589 320
rect 543 212 549 308
rect 583 212 589 308
rect 631 308 677 320
rect 631 258 637 308
rect 671 258 677 308
rect 543 200 589 212
rect 618 206 628 258
rect 680 206 690 258
rect 631 200 677 206
rect 335 172 369 200
rect 0 138 720 172
rect 323 122 382 138
rect 323 88 335 122
rect 369 88 382 122
rect 323 83 382 88
rect 323 82 381 83
<< via1 >>
rect 38 212 47 258
rect 47 212 81 258
rect 81 212 90 258
rect 38 206 90 212
rect 628 212 637 258
rect 637 212 671 258
rect 671 212 680 258
rect 628 206 680 212
<< metal2 >>
rect 38 258 90 696
rect 38 0 90 206
rect 628 258 680 696
rect 628 0 680 206
<< labels >>
rlabel metal2 628 0 680 47 0 BL_
rlabel metal1 0 138 38 172 0 VSS
rlabel metal1 0 410 22 444 0 WL
rlabel metal1 0 662 38 696 0 VDD
rlabel metal2 38 0 90 47 0 BL
<< end >>
