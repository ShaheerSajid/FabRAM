.title characterizer
.include /home/shaheer/Desktop/FabRAM/FE/out/sram256x32.spi
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

      .tran 0.011615649999999998n 23.231299999999997n 0.0n
      .control
      set hcopydevtype = svg
      run
      meas tran tdiff_cell_rise TRIG v(clk) VAL=0.9 RISE=3   TARG v(Q0) VAL=0.9 RISE=LAST 
      meas tran tdiff_tran_rise TRIG v(Q0)  VAL=0.18000000000000002 RISE=LAST TARG v(Q0) VAL=1.62 RISE=LAST 
      meas tran tdiff_cell_fall TRIG v(clk) VAL=0.9 RISE=4 TARG v(Q0) VAL=0.9 FALL=LAST 
      meas tran tdiff_tran_fall TRIG v(Q0)  VAL=1.62 FALL=LAST TARG v(Q0) VAL=0.18000000000000002 FALL=LAST 

      echo "$&tdiff_cell_rise,$&tdiff_tran_rise $&tdiff_cell_fall,$&tdiff_tran_fall" > log/sim_0.32313_0.03967.text
      hardcopy log/sim_0.32313_0.03967.svg v(clk)+10 v(x0.WLEN)+8 v(x0.DC0)+8 v(x0.WL0)+8 v(x0.DBL)+6 v(x0.DBL_)+6 v(x0.SAEN)+6 v(x0.BL0)+4 v(x0.BL_0)+4 v(x0.DR0)+2 v(x0.DR_0)+2 v(x0.DW0) v(x0.DW_0) v(Q0)-6 v(x0.WREN)-8
      exit
      .endc
      
Vpower VDD 0 1.8
Vgnd VSS 0 0
Vclk clk VSS DC 0V PULSE(0V 1.8V 0ns 0.40391249999999995ns 0.40391249999999995ns 2.5ns 5.807824999999999ns)
Vaddr addr VSS DC 0V PULSE(0V 1.8V 0s 1ps 1ps 2.5ns 11.615649999999999ns)
Vdin din VSS DC 0V PULSE(0V 1.8V 0s 1ps 1ps 2.5ns 11.615649999999999ns)
Vwrite write VSS DC 0V PULSE(0V 1.8V 0s 1ps 1ps 11.615649999999999ns 23.231299999999997ns)
X0 VDD VSS clk addr addr addr addr addr addr addr addr din din din din din din din din din din din din din din din din din din din din din din din din din din din din din din din din Q0 Q1 Q2 Q3 Q4 Q5 Q6 Q7 Q8 Q9 Q10 Q11 Q12 Q13 Q14 Q15 Q16 Q17 Q18 Q19 Q20 Q21 Q22 Q23 Q24 Q25 Q26 Q27 Q28 Q29 Q30 Q31 write VDD sram256x32
C0 Q0 VSS 0.03967p
