magic
tech sky130A
magscale 1 2
timestamp 1702544174
<< nwell >>
rect 0 1516 720 2572
rect 0 559 720 767
<< nmos >>
rect 119 1364 149 1448
rect 207 1364 237 1448
rect 467 1364 497 1448
rect 555 1364 585 1448
rect 168 970 198 1054
rect 497 970 527 1054
rect 585 970 615 1054
rect 219 117 249 317
rect 455 117 485 317
<< pmos >>
rect 293 2310 323 2510
rect 381 2310 411 2510
rect 119 2086 149 2186
rect 337 1947 367 2147
rect 555 2086 585 2186
rect 119 1578 149 1662
rect 207 1578 237 1662
rect 467 1578 497 1662
rect 555 1578 585 1662
rect 168 621 198 705
rect 497 621 527 705
rect 585 621 615 705
<< ndiff >>
rect 61 1436 119 1448
rect 61 1376 73 1436
rect 107 1376 119 1436
rect 61 1364 119 1376
rect 149 1436 207 1448
rect 149 1376 161 1436
rect 195 1376 207 1436
rect 149 1364 207 1376
rect 237 1436 295 1448
rect 237 1376 249 1436
rect 283 1376 295 1436
rect 237 1364 295 1376
rect 409 1436 467 1448
rect 409 1376 421 1436
rect 455 1376 467 1436
rect 409 1364 467 1376
rect 497 1436 555 1448
rect 497 1376 509 1436
rect 543 1376 555 1436
rect 497 1364 555 1376
rect 585 1436 643 1448
rect 585 1376 597 1436
rect 631 1376 643 1436
rect 585 1364 643 1376
rect 110 1042 168 1054
rect 110 982 122 1042
rect 156 982 168 1042
rect 110 970 168 982
rect 198 1042 256 1054
rect 198 982 210 1042
rect 244 982 256 1042
rect 198 970 256 982
rect 439 1042 497 1054
rect 439 982 451 1042
rect 485 982 497 1042
rect 439 970 497 982
rect 527 1042 585 1054
rect 527 982 539 1042
rect 573 982 585 1042
rect 527 970 585 982
rect 615 1042 673 1054
rect 615 982 627 1042
rect 661 982 673 1042
rect 615 970 673 982
rect 161 305 219 317
rect 161 129 173 305
rect 207 129 219 305
rect 161 117 219 129
rect 249 305 307 317
rect 249 129 261 305
rect 295 129 307 305
rect 249 117 307 129
rect 397 305 455 317
rect 397 129 409 305
rect 443 129 455 305
rect 397 117 455 129
rect 485 305 543 317
rect 485 129 497 305
rect 531 129 543 305
rect 485 117 543 129
<< pdiff >>
rect 235 2498 293 2510
rect 235 2322 247 2498
rect 281 2322 293 2498
rect 235 2310 293 2322
rect 323 2498 381 2510
rect 323 2322 335 2498
rect 369 2322 381 2498
rect 323 2310 381 2322
rect 411 2498 469 2510
rect 411 2322 423 2498
rect 457 2322 469 2498
rect 411 2310 469 2322
rect 61 2174 119 2186
rect 61 2098 73 2174
rect 107 2098 119 2174
rect 61 2086 119 2098
rect 149 2174 207 2186
rect 149 2098 161 2174
rect 195 2098 207 2174
rect 497 2174 555 2186
rect 149 2086 207 2098
rect 279 2135 337 2147
rect 279 1959 291 2135
rect 325 1959 337 2135
rect 279 1947 337 1959
rect 367 2135 425 2147
rect 367 1959 379 2135
rect 413 1959 425 2135
rect 497 2098 509 2174
rect 543 2098 555 2174
rect 497 2086 555 2098
rect 585 2174 643 2186
rect 585 2098 597 2174
rect 631 2098 643 2174
rect 585 2086 643 2098
rect 367 1947 425 1959
rect 61 1650 119 1662
rect 61 1590 73 1650
rect 107 1590 119 1650
rect 61 1578 119 1590
rect 149 1650 207 1662
rect 149 1590 161 1650
rect 195 1590 207 1650
rect 149 1578 207 1590
rect 237 1650 295 1662
rect 237 1590 249 1650
rect 283 1590 295 1650
rect 237 1578 295 1590
rect 409 1650 467 1662
rect 409 1590 421 1650
rect 455 1590 467 1650
rect 409 1578 467 1590
rect 497 1650 555 1662
rect 497 1590 509 1650
rect 543 1590 555 1650
rect 497 1578 555 1590
rect 585 1650 643 1662
rect 585 1590 597 1650
rect 631 1590 643 1650
rect 585 1578 643 1590
rect 110 693 168 705
rect 110 633 122 693
rect 156 633 168 693
rect 110 621 168 633
rect 198 693 256 705
rect 198 633 210 693
rect 244 633 256 693
rect 198 621 256 633
rect 439 693 497 705
rect 439 633 451 693
rect 485 633 497 693
rect 439 621 497 633
rect 527 693 585 705
rect 527 633 539 693
rect 573 633 585 693
rect 527 621 585 633
rect 615 693 673 705
rect 615 633 627 693
rect 661 633 673 693
rect 615 621 673 633
<< ndiffc >>
rect 73 1376 107 1436
rect 161 1376 195 1436
rect 249 1376 283 1436
rect 421 1376 455 1436
rect 509 1376 543 1436
rect 597 1376 631 1436
rect 122 982 156 1042
rect 210 982 244 1042
rect 451 982 485 1042
rect 539 982 573 1042
rect 627 982 661 1042
rect 173 129 207 305
rect 261 129 295 305
rect 409 129 443 305
rect 497 129 531 305
<< pdiffc >>
rect 247 2322 281 2498
rect 335 2322 369 2498
rect 423 2322 457 2498
rect 73 2098 107 2174
rect 161 2098 195 2174
rect 291 1959 325 2135
rect 379 1959 413 2135
rect 509 2098 543 2174
rect 597 2098 631 2174
rect 73 1590 107 1650
rect 161 1590 195 1650
rect 249 1590 283 1650
rect 421 1590 455 1650
rect 509 1590 543 1650
rect 597 1590 631 1650
rect 122 633 156 693
rect 210 633 244 693
rect 451 633 485 693
rect 539 633 573 693
rect 627 633 661 693
<< psubdiff >>
rect 311 1274 393 1293
rect 311 1214 335 1274
rect 369 1214 393 1274
rect 311 1185 393 1214
rect 310 1042 368 1066
rect 310 982 322 1042
rect 356 982 368 1042
rect 310 958 368 982
<< nsubdiff >>
rect 97 2387 179 2411
rect 97 2327 122 2387
rect 156 2327 179 2387
rect 97 2303 179 2327
rect 310 693 368 717
rect 310 633 322 693
rect 356 633 368 693
rect 310 609 368 633
<< psubdiffcont >>
rect 335 1214 369 1274
rect 322 982 356 1042
<< nsubdiffcont >>
rect 122 2327 156 2387
rect 322 633 356 693
<< poly >>
rect 293 2510 323 2536
rect 381 2510 411 2536
rect 293 2284 323 2310
rect 381 2284 411 2310
rect 293 2262 411 2284
rect 293 2254 334 2262
rect 318 2228 334 2254
rect 368 2254 411 2262
rect 368 2228 384 2254
rect 318 2212 384 2228
rect 119 2186 149 2212
rect 337 2147 367 2212
rect 555 2186 585 2212
rect 119 1899 149 2086
rect 337 1921 367 1947
rect 555 1899 585 2086
rect 119 1883 199 1899
rect 119 1849 135 1883
rect 169 1849 199 1883
rect 119 1833 199 1849
rect 505 1883 585 1899
rect 505 1849 535 1883
rect 569 1849 585 1883
rect 505 1833 585 1849
rect 119 1662 149 1688
rect 207 1662 237 1688
rect 467 1662 497 1688
rect 555 1662 585 1688
rect 119 1448 149 1578
rect 207 1540 237 1578
rect 207 1524 287 1540
rect 207 1490 237 1524
rect 271 1490 287 1524
rect 207 1474 287 1490
rect 207 1448 237 1474
rect 467 1448 497 1578
rect 555 1540 585 1578
rect 555 1524 635 1540
rect 555 1490 585 1524
rect 619 1490 635 1524
rect 555 1474 635 1490
rect 555 1448 585 1474
rect 119 1275 149 1364
rect 207 1338 237 1364
rect 103 1259 169 1275
rect 103 1225 119 1259
rect 153 1225 169 1259
rect 103 1209 169 1225
rect 467 1201 497 1364
rect 555 1259 585 1364
rect 555 1229 615 1259
rect 451 1185 517 1201
rect 451 1151 467 1185
rect 501 1151 517 1185
rect 451 1135 517 1151
rect 168 1054 198 1080
rect 497 1054 527 1080
rect 585 1054 615 1229
rect 168 861 198 970
rect 168 845 259 861
rect 168 811 209 845
rect 243 811 259 845
rect 168 795 259 811
rect 168 705 198 795
rect 497 705 527 970
rect 585 705 615 970
rect 168 595 198 621
rect 497 541 527 621
rect 585 595 615 621
rect 479 525 545 541
rect 479 491 495 525
rect 529 491 545 525
rect 479 475 545 491
rect 319 455 385 471
rect 319 421 335 455
rect 369 421 385 455
rect 319 415 385 421
rect 219 385 485 415
rect 219 317 249 385
rect 455 317 485 385
rect 219 91 249 117
rect 455 91 485 117
<< polycont >>
rect 334 2228 368 2262
rect 135 1849 169 1883
rect 535 1849 569 1883
rect 237 1490 271 1524
rect 585 1490 619 1524
rect 119 1225 153 1259
rect 467 1151 501 1185
rect 209 811 243 845
rect 495 491 529 525
rect 335 421 369 455
<< locali >>
rect 122 2548 369 2582
rect 122 2403 156 2548
rect 247 2498 281 2514
rect 108 2387 170 2403
rect 108 2327 122 2387
rect 156 2327 170 2387
rect 108 2311 170 2327
rect 73 2174 107 2190
rect 73 2082 107 2098
rect 161 2174 195 2190
rect 247 2156 281 2322
rect 335 2498 369 2548
rect 335 2306 369 2322
rect 423 2498 457 2514
rect 318 2228 334 2262
rect 368 2228 384 2262
rect 423 2156 457 2322
rect 247 2135 325 2156
rect 247 2122 291 2135
rect 161 1977 195 2098
rect 161 1959 291 1977
rect 161 1943 325 1959
rect 379 2135 457 2156
rect 413 2122 457 2135
rect 509 2174 543 2190
rect 509 1977 543 2098
rect 597 2174 631 2190
rect 597 2082 631 2098
rect 413 1959 543 1977
rect 379 1943 543 1959
rect 119 1849 135 1883
rect 169 1849 535 1883
rect 569 1849 632 1883
rect 195 1771 283 1805
rect 73 1650 107 1666
rect 73 1524 107 1590
rect 161 1650 195 1666
rect 161 1574 195 1590
rect 249 1650 283 1771
rect 597 1666 632 1849
rect 249 1574 283 1590
rect 421 1650 455 1666
rect 421 1524 455 1590
rect 509 1650 543 1666
rect 509 1574 543 1590
rect 597 1650 631 1666
rect 597 1574 631 1590
rect 73 1490 237 1524
rect 271 1490 287 1524
rect 421 1490 585 1524
rect 619 1490 635 1524
rect 73 1436 107 1490
rect 73 1360 107 1376
rect 161 1436 195 1452
rect 161 1360 195 1376
rect 249 1436 283 1452
rect 249 1360 283 1376
rect 421 1436 455 1490
rect 421 1360 455 1376
rect 509 1436 543 1452
rect 509 1324 543 1376
rect 597 1436 631 1452
rect 597 1360 631 1376
rect 319 1290 544 1324
rect 319 1274 385 1290
rect 103 1225 119 1259
rect 153 1225 169 1259
rect 319 1214 335 1274
rect 369 1214 385 1274
rect 319 1198 385 1214
rect 319 1058 356 1198
rect 451 1151 467 1185
rect 501 1151 517 1185
rect 122 1042 156 1058
rect 122 693 156 982
rect 210 1042 356 1058
rect 244 982 322 1042
rect 210 966 356 982
rect 451 1042 485 1058
rect 451 966 485 982
rect 539 1042 573 1058
rect 539 966 573 982
rect 627 1042 661 1058
rect 627 966 661 982
rect 193 811 209 845
rect 243 811 259 845
rect 122 455 156 633
rect 210 693 368 709
rect 244 633 322 693
rect 356 633 368 693
rect 210 617 368 633
rect 451 693 485 709
rect 451 617 485 633
rect 539 693 573 709
rect 539 617 573 633
rect 627 693 661 709
rect 627 617 661 633
rect 479 491 495 525
rect 529 491 545 525
rect 122 421 335 455
rect 369 421 385 455
rect 173 305 207 321
rect 173 113 207 129
rect 261 305 295 321
rect 261 113 295 129
rect 409 305 443 321
rect 409 113 443 129
rect 497 305 531 321
rect 497 113 531 129
<< viali >>
rect 247 2322 281 2498
rect 73 2098 107 2174
rect 161 2098 195 2174
rect 335 2322 369 2498
rect 423 2322 457 2498
rect 334 2228 368 2262
rect 291 1959 325 2135
rect 379 1959 413 2135
rect 509 2098 543 2174
rect 597 2098 631 2174
rect 161 1771 195 1805
rect 73 1590 107 1650
rect 161 1590 195 1650
rect 249 1590 283 1650
rect 421 1590 455 1650
rect 509 1590 543 1650
rect 597 1590 631 1650
rect 73 1376 107 1436
rect 161 1376 195 1436
rect 249 1376 283 1436
rect 421 1376 455 1436
rect 509 1376 543 1436
rect 597 1376 631 1436
rect 119 1225 153 1259
rect 467 1151 501 1185
rect 122 982 156 1042
rect 210 982 244 1042
rect 451 982 485 1042
rect 539 982 573 1042
rect 627 982 661 1042
rect 209 811 243 845
rect 122 633 156 693
rect 210 633 244 693
rect 451 633 485 693
rect 539 633 573 693
rect 627 633 661 693
rect 495 491 529 525
rect 173 129 207 305
rect 261 129 295 305
rect 409 129 443 305
rect 497 129 531 305
<< metal1 >>
rect 0 2556 720 2590
rect 28 2476 38 2528
rect 90 2510 100 2528
rect 335 2510 369 2556
rect 90 2498 287 2510
rect 90 2476 247 2498
rect 241 2322 247 2476
rect 281 2322 287 2498
rect 241 2310 287 2322
rect 329 2498 375 2510
rect 329 2322 335 2498
rect 369 2322 375 2498
rect 329 2310 375 2322
rect 417 2498 467 2528
rect 417 2322 423 2498
rect 457 2476 467 2498
rect 519 2476 529 2528
rect 457 2322 463 2476
rect 580 2323 614 2556
rect 417 2310 463 2322
rect 142 2222 152 2274
rect 204 2268 214 2274
rect 542 2271 552 2323
rect 604 2271 614 2323
rect 204 2262 380 2268
rect 204 2228 334 2262
rect 368 2228 384 2262
rect 204 2222 380 2228
rect 67 2174 113 2186
rect 67 2098 73 2174
rect 107 2098 113 2174
rect 67 2086 113 2098
rect 155 2174 201 2186
rect 155 2098 161 2174
rect 195 2098 201 2174
rect 503 2174 549 2186
rect 155 2086 201 2098
rect 285 2135 331 2147
rect 54 2034 64 2086
rect 116 2034 126 2086
rect 285 1999 291 2135
rect 242 1947 252 1999
rect 325 1959 331 2135
rect 304 1947 331 1959
rect 373 2135 419 2147
rect 373 1959 379 2135
rect 413 1999 419 2135
rect 503 2098 509 2174
rect 543 2098 549 2174
rect 503 2086 549 2098
rect 591 2174 637 2186
rect 591 2098 597 2174
rect 631 2098 637 2174
rect 591 2086 637 2098
rect 578 2034 588 2086
rect 640 2034 650 2086
rect 373 1947 400 1959
rect 452 1947 462 1999
rect 142 1762 152 1814
rect 204 1762 214 1814
rect 490 1734 500 1752
rect 0 1700 500 1734
rect 552 1734 562 1752
rect 552 1700 720 1734
rect 161 1662 195 1700
rect 67 1650 113 1662
rect 67 1590 73 1650
rect 107 1590 113 1650
rect 67 1578 113 1590
rect 155 1650 201 1662
rect 155 1590 161 1650
rect 195 1590 201 1650
rect 155 1578 201 1590
rect 243 1650 289 1662
rect 243 1590 249 1650
rect 283 1590 289 1650
rect 243 1578 289 1590
rect 249 1448 283 1578
rect 335 1526 369 1700
rect 509 1662 543 1700
rect 415 1650 461 1662
rect 415 1590 421 1650
rect 455 1590 461 1650
rect 415 1578 461 1590
rect 503 1650 549 1662
rect 503 1590 509 1650
rect 543 1590 549 1650
rect 503 1578 549 1590
rect 591 1650 637 1662
rect 591 1590 597 1650
rect 631 1590 637 1650
rect 591 1578 637 1590
rect 316 1474 326 1526
rect 378 1474 388 1526
rect 597 1448 631 1578
rect 67 1436 113 1448
rect 67 1376 73 1436
rect 107 1376 113 1436
rect 67 1364 113 1376
rect 155 1436 201 1448
rect 155 1376 161 1436
rect 195 1376 201 1436
rect 155 1364 201 1376
rect 243 1436 289 1448
rect 243 1376 249 1436
rect 283 1376 289 1436
rect 243 1364 289 1376
rect 415 1436 461 1448
rect 415 1376 421 1436
rect 455 1376 461 1436
rect 415 1364 461 1376
rect 503 1436 549 1448
rect 503 1376 509 1436
rect 543 1376 549 1436
rect 503 1364 549 1376
rect 591 1436 637 1448
rect 591 1376 597 1436
rect 631 1376 637 1436
rect 591 1364 637 1376
rect 161 1327 195 1364
rect 509 1327 543 1364
rect 0 1293 720 1327
rect 107 1259 165 1265
rect 0 1225 119 1259
rect 153 1225 720 1259
rect 107 1219 165 1225
rect 516 1191 526 1197
rect 455 1185 526 1191
rect 455 1151 467 1185
rect 501 1151 526 1185
rect 455 1145 526 1151
rect 578 1145 588 1197
rect 0 1083 720 1117
rect 210 1054 244 1083
rect 451 1054 485 1083
rect 627 1054 661 1083
rect 116 1042 162 1054
rect 116 982 122 1042
rect 156 982 162 1042
rect 116 970 162 982
rect 204 1042 250 1054
rect 204 982 210 1042
rect 244 982 250 1042
rect 204 970 250 982
rect 445 1042 491 1054
rect 445 982 451 1042
rect 485 982 491 1042
rect 445 970 491 982
rect 533 1042 579 1054
rect 533 982 539 1042
rect 573 982 579 1042
rect 533 970 579 982
rect 621 1042 667 1054
rect 621 982 627 1042
rect 661 982 667 1042
rect 621 970 667 982
rect 197 845 255 851
rect 539 845 573 970
rect 197 811 209 845
rect 243 811 573 845
rect 197 805 255 811
rect 539 705 573 811
rect 116 693 162 705
rect 116 633 122 693
rect 156 633 162 693
rect 116 621 162 633
rect 204 693 250 705
rect 204 633 210 693
rect 244 633 250 693
rect 445 693 491 705
rect 204 621 250 633
rect 210 593 244 621
rect 316 593 326 645
rect 378 593 388 645
rect 445 633 451 693
rect 485 633 491 693
rect 445 621 491 633
rect 533 693 579 705
rect 533 633 539 693
rect 573 633 579 693
rect 533 621 579 633
rect 621 693 667 705
rect 621 633 627 693
rect 661 633 667 693
rect 621 621 667 633
rect 451 593 485 621
rect 627 593 661 621
rect 0 559 720 593
rect 483 525 541 531
rect 0 491 495 525
rect 529 491 720 525
rect 483 485 541 491
rect 316 411 326 463
rect 378 455 388 463
rect 378 421 588 455
rect 378 411 388 421
rect 516 369 526 421
rect 578 369 588 421
rect 242 317 252 369
rect 304 317 314 369
rect 390 317 400 369
rect 452 317 462 369
rect 167 305 213 317
rect 167 129 173 305
rect 207 129 213 305
rect 167 117 213 129
rect 255 305 301 317
rect 255 129 261 305
rect 295 129 301 305
rect 255 117 301 129
rect 403 305 449 317
rect 403 129 409 305
rect 443 129 449 305
rect 403 117 449 129
rect 491 305 537 317
rect 491 129 497 305
rect 531 129 537 305
rect 491 117 537 129
rect 154 65 164 117
rect 216 65 226 117
rect 478 65 488 117
rect 540 65 550 117
<< via1 >>
rect 38 2476 90 2528
rect 467 2476 519 2528
rect 152 2222 204 2274
rect 552 2271 604 2323
rect 64 2034 116 2086
rect 252 1959 291 1999
rect 291 1959 304 1999
rect 252 1947 304 1959
rect 588 2034 640 2086
rect 400 1959 413 1999
rect 413 1959 452 1999
rect 400 1947 452 1959
rect 152 1805 204 1814
rect 152 1771 161 1805
rect 161 1771 195 1805
rect 195 1771 204 1805
rect 152 1762 204 1771
rect 500 1700 552 1752
rect 326 1474 378 1526
rect 526 1145 578 1197
rect 326 593 378 645
rect 326 411 378 463
rect 526 369 578 421
rect 252 317 304 369
rect 400 317 452 369
rect 164 65 216 117
rect 488 65 540 117
<< metal2 >>
rect 38 2528 90 2624
rect 38 2466 90 2476
rect 467 2528 519 2538
rect 628 2528 680 2624
rect 519 2476 680 2528
rect 467 2466 519 2476
rect 500 2323 604 2333
rect 152 2274 204 2284
rect 64 2086 116 2096
rect 64 1263 116 2034
rect 152 1814 204 2222
rect 500 2271 552 2323
rect 500 2261 604 2271
rect 152 1752 204 1762
rect 252 1999 304 2009
rect 252 1616 304 1947
rect 12 1235 116 1263
rect 207 1564 304 1616
rect 400 1999 452 2009
rect 400 1616 452 1947
rect 500 1752 552 2261
rect 500 1690 552 1700
rect 588 2086 640 2096
rect 400 1564 497 1616
rect 12 0 64 1235
rect 207 377 259 1564
rect 326 1526 378 1536
rect 326 645 378 1474
rect 326 583 378 593
rect 326 463 378 473
rect 326 405 378 411
rect 207 369 304 377
rect 207 317 252 369
rect 207 309 304 317
rect 332 195 372 405
rect 445 377 497 1564
rect 588 1263 640 2034
rect 588 1235 692 1263
rect 400 369 497 377
rect 452 317 497 369
rect 526 1197 578 1207
rect 526 421 578 1145
rect 526 359 578 369
rect 400 310 497 317
rect 164 117 216 127
rect 164 0 216 65
rect 326 0 378 195
rect 488 117 540 126
rect 488 0 540 65
rect 640 0 692 1235
<< labels >>
rlabel metal1 1 491 35 525 0 WREN
rlabel metal1 1 559 35 593 0 VDD
rlabel metal1 1 1083 35 1117 0 VSS
rlabel metal1 1 1225 35 1259 0 PCHG
rlabel metal1 1 1293 35 1327 0 VSS
rlabel metal1 0 1700 34 1734 0 VDD
rlabel metal2 640 0 692 52 0 DR_
rlabel metal2 488 0 540 52 0 DW_
rlabel metal2 326 0 378 52 0 SEL
rlabel metal2 164 0 216 52 0 DW
rlabel metal2 12 0 64 52 0 DR
rlabel metal2 628 2572 680 2624 0 BL_
rlabel metal2 38 2572 90 2624 0 BL
<< end >>
