magic
tech sky130A
magscale 1 2
timestamp 1702719154
<< nwell >>
rect 0 350 2686 558
<< nmos >>
rect 197 63 227 147
rect 285 63 315 147
rect 614 63 644 147
rect 702 63 732 147
rect 920 63 950 147
rect 1198 73 1228 157
rect 1286 73 1316 157
rect 1504 72 1534 156
rect 1812 70 1842 154
rect 2126 72 2156 156
rect 2214 72 2244 156
rect 2432 72 2462 156
<< pmos >>
rect 197 412 227 496
rect 285 412 315 496
rect 614 412 644 496
rect 702 412 732 496
rect 920 412 950 496
rect 1198 412 1228 496
rect 1286 412 1316 496
rect 1504 412 1534 496
rect 1812 412 1842 496
rect 2126 412 2156 496
rect 2214 412 2244 496
rect 2432 412 2462 496
<< ndiff >>
rect 139 135 197 147
rect 139 75 151 135
rect 185 75 197 135
rect 139 63 197 75
rect 227 135 285 147
rect 227 75 239 135
rect 273 75 285 135
rect 227 63 285 75
rect 315 135 373 147
rect 315 75 327 135
rect 361 75 373 135
rect 315 63 373 75
rect 556 135 614 147
rect 556 75 568 135
rect 602 75 614 135
rect 556 63 614 75
rect 644 135 702 147
rect 644 75 656 135
rect 690 75 702 135
rect 644 63 702 75
rect 732 135 790 147
rect 732 75 744 135
rect 778 75 790 135
rect 732 63 790 75
rect 862 135 920 147
rect 862 75 874 135
rect 908 75 920 135
rect 862 63 920 75
rect 950 135 1008 147
rect 950 75 962 135
rect 996 75 1008 135
rect 950 63 1008 75
rect 1140 145 1198 157
rect 1140 85 1152 145
rect 1186 85 1198 145
rect 1140 73 1198 85
rect 1228 145 1286 157
rect 1228 85 1240 145
rect 1274 85 1286 145
rect 1228 73 1286 85
rect 1316 145 1374 157
rect 1316 85 1328 145
rect 1362 85 1374 145
rect 1316 73 1374 85
rect 1446 144 1504 156
rect 1446 84 1458 144
rect 1492 84 1504 144
rect 1446 72 1504 84
rect 1534 144 1592 156
rect 1534 84 1546 144
rect 1580 84 1592 144
rect 1534 72 1592 84
rect 1754 142 1812 154
rect 1754 82 1766 142
rect 1800 82 1812 142
rect 1754 70 1812 82
rect 1842 142 1900 154
rect 1842 82 1854 142
rect 1888 82 1900 142
rect 1842 70 1900 82
rect 2068 144 2126 156
rect 2068 84 2080 144
rect 2114 84 2126 144
rect 2068 72 2126 84
rect 2156 144 2214 156
rect 2156 84 2168 144
rect 2202 84 2214 144
rect 2156 72 2214 84
rect 2244 144 2302 156
rect 2244 84 2256 144
rect 2290 84 2302 144
rect 2244 72 2302 84
rect 2374 144 2432 156
rect 2374 84 2386 144
rect 2420 84 2432 144
rect 2374 72 2432 84
rect 2462 144 2520 156
rect 2462 84 2474 144
rect 2508 84 2520 144
rect 2462 72 2520 84
<< pdiff >>
rect 139 484 197 496
rect 139 424 151 484
rect 185 424 197 484
rect 139 412 197 424
rect 227 484 285 496
rect 227 424 239 484
rect 273 424 285 484
rect 227 412 285 424
rect 315 484 373 496
rect 315 424 327 484
rect 361 424 373 484
rect 315 412 373 424
rect 556 484 614 496
rect 556 424 568 484
rect 602 424 614 484
rect 556 412 614 424
rect 644 484 702 496
rect 644 424 656 484
rect 690 424 702 484
rect 644 412 702 424
rect 732 484 790 496
rect 732 424 744 484
rect 778 424 790 484
rect 732 412 790 424
rect 862 484 920 496
rect 862 424 874 484
rect 908 424 920 484
rect 862 412 920 424
rect 950 484 1008 496
rect 950 424 962 484
rect 996 424 1008 484
rect 950 412 1008 424
rect 1140 484 1198 496
rect 1140 424 1152 484
rect 1186 424 1198 484
rect 1140 412 1198 424
rect 1228 484 1286 496
rect 1228 424 1240 484
rect 1274 424 1286 484
rect 1228 412 1286 424
rect 1316 484 1374 496
rect 1316 424 1328 484
rect 1362 424 1374 484
rect 1316 412 1374 424
rect 1446 484 1504 496
rect 1446 424 1458 484
rect 1492 424 1504 484
rect 1446 412 1504 424
rect 1534 484 1592 496
rect 1534 424 1546 484
rect 1580 424 1592 484
rect 1534 412 1592 424
rect 1754 484 1812 496
rect 1754 424 1766 484
rect 1800 424 1812 484
rect 1754 412 1812 424
rect 1842 484 1900 496
rect 1842 424 1854 484
rect 1888 424 1900 484
rect 1842 412 1900 424
rect 2068 484 2126 496
rect 2068 424 2080 484
rect 2114 424 2126 484
rect 2068 412 2126 424
rect 2156 484 2214 496
rect 2156 424 2168 484
rect 2202 424 2214 484
rect 2156 412 2214 424
rect 2244 484 2302 496
rect 2244 424 2256 484
rect 2290 424 2302 484
rect 2244 412 2302 424
rect 2374 484 2432 496
rect 2374 424 2386 484
rect 2420 424 2432 484
rect 2374 412 2432 424
rect 2462 484 2520 496
rect 2462 424 2474 484
rect 2508 424 2520 484
rect 2462 412 2520 424
<< ndiffc >>
rect 151 75 185 135
rect 239 75 273 135
rect 327 75 361 135
rect 568 75 602 135
rect 656 75 690 135
rect 744 75 778 135
rect 874 75 908 135
rect 962 75 996 135
rect 1152 85 1186 145
rect 1240 85 1274 145
rect 1328 85 1362 145
rect 1458 84 1492 144
rect 1546 84 1580 144
rect 1766 82 1800 142
rect 1854 82 1888 142
rect 2080 84 2114 144
rect 2168 84 2202 144
rect 2256 84 2290 144
rect 2386 84 2420 144
rect 2474 84 2508 144
<< pdiffc >>
rect 151 424 185 484
rect 239 424 273 484
rect 327 424 361 484
rect 568 424 602 484
rect 656 424 690 484
rect 744 424 778 484
rect 874 424 908 484
rect 962 424 996 484
rect 1152 424 1186 484
rect 1240 424 1274 484
rect 1328 424 1362 484
rect 1458 424 1492 484
rect 1546 424 1580 484
rect 1766 424 1800 484
rect 1854 424 1888 484
rect 2080 424 2114 484
rect 2168 424 2202 484
rect 2256 424 2290 484
rect 2386 424 2420 484
rect 2474 424 2508 484
<< psubdiff >>
rect 427 114 485 138
rect 427 54 439 114
rect 473 54 485 114
rect 427 30 485 54
<< nsubdiff >>
rect 442 484 500 508
rect 442 424 454 484
rect 488 424 500 484
rect 442 400 500 424
<< psubdiffcont >>
rect 439 54 473 114
<< nsubdiffcont >>
rect 454 424 488 484
<< poly >>
rect 197 496 227 522
rect 285 496 315 522
rect 614 496 644 522
rect 702 496 732 522
rect 920 496 950 522
rect 1198 496 1228 522
rect 1286 496 1316 522
rect 1504 496 1534 522
rect 1812 496 1842 522
rect 2126 496 2156 522
rect 2214 496 2244 522
rect 2432 496 2462 522
rect 51 350 111 366
rect 197 350 227 412
rect 51 316 67 350
rect 101 316 227 350
rect 51 300 111 316
rect 197 147 227 316
rect 285 366 315 412
rect 285 350 365 366
rect 285 316 315 350
rect 349 316 365 350
rect 285 300 365 316
rect 285 147 315 300
rect 467 219 533 235
rect 614 219 644 412
rect 467 185 483 219
rect 517 185 644 219
rect 467 169 533 185
rect 614 147 644 185
rect 702 235 732 412
rect 920 374 950 412
rect 920 358 1000 374
rect 920 324 950 358
rect 984 324 1000 358
rect 920 308 1000 324
rect 1046 297 1112 313
rect 1198 297 1228 412
rect 1046 263 1062 297
rect 1096 263 1228 297
rect 920 236 1001 252
rect 1046 247 1112 263
rect 702 219 782 235
rect 702 185 732 219
rect 766 185 782 219
rect 702 169 782 185
rect 920 202 950 236
rect 984 202 1001 236
rect 920 185 1001 202
rect 702 147 732 169
rect 920 147 950 185
rect 1198 157 1228 263
rect 1286 364 1316 412
rect 1504 364 1534 412
rect 1812 364 1842 412
rect 1286 348 1366 364
rect 1286 314 1316 348
rect 1350 314 1366 348
rect 1286 298 1366 314
rect 1504 348 1584 364
rect 1504 314 1534 348
rect 1568 314 1584 348
rect 1504 298 1584 314
rect 1812 348 1892 364
rect 1812 314 1842 348
rect 1876 314 1892 348
rect 1812 298 1892 314
rect 1976 335 2042 351
rect 2126 335 2156 412
rect 1976 300 1992 335
rect 2026 300 2156 335
rect 1286 157 1316 298
rect 1976 284 2042 300
rect 1600 222 1666 238
rect 1600 202 1616 222
rect 1504 188 1616 202
rect 1650 188 1666 222
rect 1908 222 1974 238
rect 1908 210 1924 222
rect 1504 172 1666 188
rect 1812 188 1924 210
rect 1958 188 1974 222
rect 1812 180 1974 188
rect 197 37 227 63
rect 285 37 315 63
rect 1504 156 1534 172
rect 614 37 644 63
rect 702 37 732 63
rect 920 37 950 63
rect 1198 47 1228 73
rect 1286 47 1316 73
rect 1812 154 1842 180
rect 1908 172 1974 180
rect 2126 156 2156 300
rect 2214 351 2244 412
rect 2432 374 2462 412
rect 2432 358 2512 374
rect 2214 335 2294 351
rect 2214 300 2244 335
rect 2278 300 2294 335
rect 2432 324 2462 358
rect 2496 324 2512 358
rect 2432 308 2512 324
rect 2214 284 2294 300
rect 2214 156 2244 284
rect 2432 246 2512 262
rect 2432 212 2462 246
rect 2496 212 2512 246
rect 2432 196 2512 212
rect 2432 156 2462 196
rect 1504 46 1534 72
rect 1812 44 1842 70
rect 2126 46 2156 72
rect 2214 46 2244 72
rect 2432 46 2462 72
<< polycont >>
rect 67 316 101 350
rect 315 316 349 350
rect 483 185 517 219
rect 950 324 984 358
rect 1062 263 1096 297
rect 732 185 766 219
rect 950 202 984 236
rect 1316 314 1350 348
rect 1534 314 1568 348
rect 1842 314 1876 348
rect 1992 300 2026 335
rect 1616 188 1650 222
rect 1924 188 1958 222
rect 2244 300 2278 335
rect 2462 324 2496 358
rect 2462 212 2496 246
<< locali >>
rect 151 484 185 500
rect 151 350 185 424
rect 239 484 273 500
rect 239 408 273 424
rect 327 484 361 500
rect 327 408 361 424
rect 454 484 488 500
rect 454 408 488 424
rect 568 484 602 500
rect 51 316 67 350
rect 101 316 117 350
rect 151 316 315 350
rect 349 316 447 350
rect 151 135 185 316
rect 413 297 447 316
rect 568 219 602 424
rect 656 484 690 500
rect 656 408 690 424
rect 744 484 778 500
rect 874 484 908 500
rect 778 438 874 472
rect 744 408 778 424
rect 273 185 483 219
rect 517 185 533 219
rect 568 185 732 219
rect 766 185 782 219
rect 151 59 185 75
rect 239 135 273 151
rect 239 59 273 75
rect 327 135 361 151
rect 568 135 602 185
rect 327 59 361 75
rect 439 114 473 130
rect 568 59 602 75
rect 656 135 690 151
rect 656 59 690 75
rect 744 135 778 151
rect 874 135 908 424
rect 962 484 996 500
rect 1152 484 1186 500
rect 996 424 1096 442
rect 962 408 1096 424
rect 950 358 984 374
rect 950 308 984 324
rect 1062 297 1096 408
rect 950 236 984 252
rect 950 185 984 202
rect 1062 151 1096 263
rect 778 89 874 123
rect 744 59 778 75
rect 874 59 908 75
rect 962 135 1096 151
rect 996 117 1096 135
rect 1152 348 1186 424
rect 1240 484 1274 500
rect 1240 408 1274 424
rect 1328 484 1362 500
rect 1458 484 1492 500
rect 1362 438 1458 472
rect 1328 408 1362 424
rect 1152 314 1316 348
rect 1350 314 1366 348
rect 1152 145 1186 314
rect 962 59 996 75
rect 439 38 473 54
rect 1152 34 1186 85
rect 1240 145 1274 161
rect 1240 69 1274 85
rect 1328 145 1362 161
rect 1458 144 1492 424
rect 1546 484 1580 500
rect 1766 484 1800 500
rect 1580 438 1718 472
rect 1546 408 1580 424
rect 1534 348 1568 364
rect 1534 228 1568 314
rect 1616 222 1650 350
rect 1616 172 1650 188
rect 1684 297 1718 438
rect 1362 89 1458 123
rect 1328 69 1362 85
rect 1458 68 1492 84
rect 1546 144 1580 160
rect 1684 120 1718 263
rect 1580 86 1718 120
rect 1766 142 1800 424
rect 1854 484 1888 500
rect 2080 484 2114 500
rect 1888 438 2026 472
rect 1854 408 1888 424
rect 1842 348 1876 364
rect 1842 227 1876 314
rect 1924 222 1958 350
rect 1924 172 1958 188
rect 1992 335 2026 438
rect 1546 68 1580 84
rect 1766 34 1800 82
rect 1854 142 1888 158
rect 1992 120 2026 300
rect 1888 86 2026 120
rect 1854 66 1888 82
rect 1152 0 1800 34
rect 1992 34 2026 86
rect 2080 335 2114 424
rect 2168 484 2202 500
rect 2168 408 2202 424
rect 2256 484 2290 500
rect 2386 484 2420 500
rect 2290 437 2386 471
rect 2256 408 2290 424
rect 2080 301 2244 335
rect 2114 300 2244 301
rect 2278 300 2294 335
rect 2080 144 2114 267
rect 2080 68 2114 84
rect 2168 144 2202 160
rect 2168 68 2202 84
rect 2256 144 2290 160
rect 2386 144 2420 424
rect 2474 484 2508 500
rect 2508 424 2569 442
rect 2474 408 2569 424
rect 2462 358 2496 374
rect 2462 308 2496 324
rect 2462 246 2496 262
rect 2462 196 2496 212
rect 2535 160 2569 408
rect 2290 96 2386 130
rect 2256 68 2290 84
rect 2386 68 2420 84
rect 2474 144 2569 160
rect 2508 125 2569 144
rect 2474 34 2508 84
rect 1992 0 2508 34
<< viali >>
rect 151 424 185 484
rect 239 424 273 484
rect 327 424 361 484
rect 454 437 488 471
rect 568 424 602 484
rect 67 316 101 350
rect 413 263 447 297
rect 656 424 690 484
rect 744 424 778 484
rect 874 424 908 484
rect 239 185 273 219
rect 151 75 185 135
rect 239 75 273 135
rect 327 75 361 135
rect 439 67 473 101
rect 568 75 602 135
rect 656 75 690 135
rect 744 75 778 135
rect 962 424 996 484
rect 950 324 984 358
rect 1062 263 1096 297
rect 950 202 984 236
rect 874 75 908 135
rect 962 75 996 135
rect 1152 424 1186 484
rect 1240 424 1274 484
rect 1328 424 1362 484
rect 1458 424 1492 484
rect 1152 85 1186 145
rect 1240 85 1274 145
rect 1328 85 1362 145
rect 1546 424 1580 484
rect 1534 194 1568 228
rect 1616 350 1650 384
rect 1684 263 1718 297
rect 1458 84 1492 144
rect 1546 84 1580 144
rect 1766 424 1800 484
rect 1854 424 1888 484
rect 1842 193 1876 227
rect 1924 350 1958 384
rect 1766 82 1800 142
rect 1854 82 1888 142
rect 2080 424 2114 484
rect 2168 424 2202 484
rect 2256 424 2290 484
rect 2386 424 2420 484
rect 2080 267 2114 301
rect 2080 84 2114 144
rect 2168 84 2202 144
rect 2256 84 2290 144
rect 2474 424 2508 484
rect 2462 324 2496 358
rect 2462 212 2496 246
rect 2386 84 2420 144
rect 2474 84 2508 144
<< metal1 >>
rect 0 524 2686 558
rect 239 496 273 524
rect 145 484 191 496
rect 145 424 151 484
rect 185 424 191 484
rect 145 412 191 424
rect 233 484 279 496
rect 233 424 239 484
rect 273 424 279 484
rect 233 412 279 424
rect 321 484 367 496
rect 321 424 327 484
rect 361 424 367 484
rect 454 477 488 524
rect 656 496 690 524
rect 1240 496 1274 524
rect 2168 496 2202 524
rect 562 484 608 496
rect 442 471 500 477
rect 442 437 454 471
rect 488 437 500 471
rect 442 431 500 437
rect 321 412 367 424
rect 562 424 568 484
rect 602 424 608 484
rect 562 412 608 424
rect 650 484 696 496
rect 650 424 656 484
rect 690 424 696 484
rect 650 412 696 424
rect 738 484 784 496
rect 738 424 744 484
rect 778 424 784 484
rect 738 412 784 424
rect 868 484 914 496
rect 868 424 874 484
rect 908 424 914 484
rect 868 412 914 424
rect 956 484 1002 496
rect 956 424 962 484
rect 996 424 1002 484
rect 956 412 1002 424
rect 1146 484 1192 496
rect 1146 424 1152 484
rect 1186 424 1192 484
rect 1146 412 1192 424
rect 1234 484 1280 496
rect 1234 424 1240 484
rect 1274 424 1280 484
rect 1234 412 1280 424
rect 1322 484 1368 496
rect 1322 424 1328 484
rect 1362 424 1368 484
rect 1322 412 1368 424
rect 1452 484 1498 496
rect 1452 424 1458 484
rect 1492 424 1498 484
rect 1452 412 1498 424
rect 1540 484 1586 496
rect 1540 424 1546 484
rect 1580 424 1586 484
rect 1540 412 1586 424
rect 1760 484 1806 496
rect 1760 424 1766 484
rect 1800 424 1806 484
rect 1760 412 1806 424
rect 1848 484 1894 496
rect 1848 424 1854 484
rect 1888 424 1894 484
rect 1848 412 1894 424
rect 2074 484 2120 496
rect 2074 424 2080 484
rect 2114 424 2120 484
rect 2074 412 2120 424
rect 2162 484 2208 496
rect 2162 424 2168 484
rect 2202 424 2208 484
rect 2162 412 2208 424
rect 2250 484 2296 496
rect 2250 424 2256 484
rect 2290 424 2296 484
rect 2250 412 2296 424
rect 2380 484 2426 496
rect 2380 424 2386 484
rect 2420 424 2426 484
rect 2380 412 2426 424
rect 2468 484 2514 496
rect 2468 424 2474 484
rect 2508 424 2514 484
rect 2468 412 2514 424
rect 327 384 361 412
rect 1604 384 1662 390
rect 1912 384 1970 390
rect 327 358 1616 384
rect 55 350 113 356
rect 0 316 67 350
rect 101 316 113 350
rect 55 310 113 316
rect 327 350 950 358
rect 227 219 285 225
rect 0 185 239 219
rect 273 185 285 219
rect 227 179 285 185
rect 327 147 361 350
rect 938 324 950 350
rect 984 350 1616 358
rect 1650 350 1924 384
rect 1958 358 2508 384
rect 1958 350 2462 358
rect 984 324 996 350
rect 1604 344 1662 350
rect 1912 344 1970 350
rect 938 318 996 324
rect 2450 324 2462 350
rect 2496 324 2508 358
rect 2450 318 2508 324
rect 401 297 459 303
rect 401 263 413 297
rect 447 263 459 297
rect 401 257 459 263
rect 1050 297 1108 303
rect 1672 297 1730 303
rect 1050 263 1062 297
rect 1096 263 1684 297
rect 1718 263 1730 297
rect 1050 257 1108 263
rect 1672 257 1730 263
rect 2061 258 2071 310
rect 2123 258 2133 310
rect 2559 262 2569 314
rect 2621 306 2631 314
rect 2621 272 2686 306
rect 2621 262 2631 272
rect 413 219 447 257
rect 2449 246 2508 254
rect 938 236 996 242
rect 938 219 950 236
rect 413 202 950 219
rect 984 219 996 236
rect 1522 228 1580 234
rect 1522 219 1534 228
rect 984 202 1534 219
rect 413 194 1534 202
rect 1568 219 1580 228
rect 1830 227 1888 233
rect 1830 219 1842 227
rect 1568 194 1842 219
rect 413 193 1842 194
rect 1876 219 1888 227
rect 2449 219 2462 246
rect 1876 212 2462 219
rect 2496 212 2508 246
rect 1876 193 2508 212
rect 413 185 2508 193
rect 145 135 191 147
rect 145 75 151 135
rect 185 75 191 135
rect 145 63 191 75
rect 233 135 279 147
rect 233 75 239 135
rect 273 75 279 135
rect 233 63 279 75
rect 321 135 367 147
rect 321 75 327 135
rect 361 75 367 135
rect 562 135 608 147
rect 321 63 367 75
rect 427 101 485 107
rect 427 67 439 101
rect 473 67 485 101
rect 239 34 273 63
rect 427 34 485 67
rect 562 75 568 135
rect 602 75 608 135
rect 562 63 608 75
rect 650 135 696 147
rect 650 75 656 135
rect 690 75 696 135
rect 650 63 696 75
rect 738 135 784 147
rect 738 75 744 135
rect 778 75 784 135
rect 738 63 784 75
rect 868 135 914 147
rect 868 75 874 135
rect 908 75 914 135
rect 868 63 914 75
rect 956 135 1002 147
rect 956 75 962 135
rect 996 75 1002 135
rect 956 63 1002 75
rect 1146 145 1192 157
rect 1146 85 1152 145
rect 1186 85 1192 145
rect 1146 73 1192 85
rect 1234 145 1280 157
rect 1234 85 1240 145
rect 1274 85 1280 145
rect 1234 73 1280 85
rect 1322 145 1368 157
rect 1322 85 1328 145
rect 1362 85 1368 145
rect 1322 73 1368 85
rect 1452 144 1498 156
rect 1452 84 1458 144
rect 1492 84 1498 144
rect 656 34 690 63
rect 1240 34 1274 73
rect 1452 72 1498 84
rect 1540 144 1586 156
rect 1540 84 1546 144
rect 1580 84 1586 144
rect 1540 72 1586 84
rect 1760 142 1806 154
rect 1760 82 1766 142
rect 1800 82 1806 142
rect 1760 70 1806 82
rect 1848 142 1894 154
rect 1848 82 1854 142
rect 1888 82 1894 142
rect 1848 70 1894 82
rect 2074 144 2120 156
rect 2074 84 2080 144
rect 2114 84 2120 144
rect 2074 72 2120 84
rect 2162 144 2208 156
rect 2162 84 2168 144
rect 2202 84 2208 144
rect 2162 72 2208 84
rect 2250 144 2296 156
rect 2250 84 2256 144
rect 2290 84 2296 144
rect 2250 72 2296 84
rect 2380 144 2426 156
rect 2380 84 2386 144
rect 2420 84 2426 144
rect 2380 72 2426 84
rect 2468 144 2514 156
rect 2468 84 2474 144
rect 2508 84 2514 144
rect 2468 72 2514 84
rect 2168 34 2202 72
rect 0 33 1274 34
rect 1921 33 2364 34
rect 0 0 2686 33
<< via1 >>
rect 2071 301 2123 310
rect 2071 267 2080 301
rect 2080 267 2114 301
rect 2114 267 2123 301
rect 2071 258 2123 267
rect 2569 262 2621 314
<< metal2 >>
rect 2071 310 2123 320
rect 2569 314 2621 324
rect 2123 271 2569 305
rect 2071 248 2123 258
rect 2569 252 2621 262
<< labels >>
rlabel metal1 0 316 34 350 0 clk
rlabel metal1 0 185 34 219 0 d
rlabel metal1 0 524 34 558 0 VDD
rlabel metal1 0 0 34 34 0 VSS
rlabel metal1 2652 272 2686 306 0 q
<< end >>
