magic
tech sky130A
magscale 1 2
timestamp 1702731179
<< poly >>
rect 94 3174 124 3252
rect 193 3230 260 3247
rect 312 3230 342 3252
rect 193 3195 209 3230
rect 243 3195 342 3230
rect 193 3179 260 3195
rect 312 3174 342 3195
rect 94 2702 124 2722
rect 94 2686 174 2702
rect 94 2652 124 2686
rect 158 2652 174 2686
rect 94 2636 174 2652
<< polycont >>
rect 209 3195 243 3230
rect 124 2652 158 2686
<< locali >>
rect 136 3230 170 3274
rect 136 3195 209 3230
rect 243 3195 260 3230
rect 136 3152 170 3195
rect 108 2652 124 2686
rect 158 2652 174 2686
<< viali >>
rect 124 2652 158 2686
<< metal1 >>
rect 466 3861 500 3901
rect 466 3827 612 3861
rect 48 3758 469 3792
rect 48 3678 82 3758
rect 117 3678 127 3730
rect 179 3678 189 3730
rect 266 3678 300 3758
rect 335 3678 345 3730
rect 397 3678 407 3730
rect 47 3176 301 3210
rect 47 3148 82 3176
rect 266 3148 301 3176
rect 354 3136 388 3290
rect 435 3225 469 3758
rect 578 3566 612 3827
rect 568 3514 578 3566
rect 630 3514 640 3566
rect 435 3191 559 3225
rect 47 2720 82 2748
rect 0 2686 82 2720
rect 112 2686 170 2692
rect 525 2686 559 3191
rect 112 2652 124 2686
rect 158 2652 286 2686
rect 112 2646 170 2652
rect 244 2631 252 2652
rect 620 85 630 137
rect 682 85 692 137
rect 620 0 654 85
<< via1 >>
rect 127 3678 179 3730
rect 345 3678 397 3730
rect 578 3514 630 3566
rect 630 85 682 137
<< metal2 >>
rect 167 3740 219 3901
rect 127 3730 219 3740
rect 179 3678 219 3730
rect 127 3668 219 3678
rect 345 3730 397 3740
rect 491 3730 543 3901
rect 397 3678 543 3730
rect 345 3668 397 3678
rect 578 3566 630 3576
rect 578 147 630 3514
rect 578 137 682 147
rect 578 85 630 137
rect 630 75 682 85
use sky130_fd_pr__nfet_01v8_JB3UY8  m1
timestamp 1702731179
transform 1 0 109 0 1 3478
box -73 -226 73 226
use sky130_fd_pr__pfet_01v8_5YUHNA  m2
timestamp 1702731179
transform 1 0 109 0 1 2948
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_5YUHNA  m3
timestamp 1702731179
transform 1 0 327 0 1 2948
box -109 -262 109 262
use sky130_fd_pr__nfet_01v8_JB3UY8  m4
timestamp 1702731179
transform 1 0 327 0 1 3478
box -73 -226 73 226
use ms_ff_f  ms_ff_f_0 ~/Desktop/FabRAM/FE/sram130/ms_ff
timestamp 1702719154
transform 0 -1 558 1 0 0
box 0 0 2686 558
<< end >>
