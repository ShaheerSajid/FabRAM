magic
tech sky130A
magscale 1 2
timestamp 1702540635
<< nwell >>
rect -199 0 0 324
rect 306 290 521 324
rect 258 218 521 290
rect 19 0 262 1
rect 306 0 521 218
rect -199 -224 -174 0
rect 44 -39 262 0
rect 44 -208 46 -39
rect 480 -224 521 0
rect -199 -524 521 -224
rect -199 -732 -174 -524
rect 132 -732 174 -524
rect 480 -732 521 -524
rect -198 -1689 -125 -1481
rect 510 -1689 522 -1481
<< psubdiff >>
rect 112 -974 194 -955
rect 112 -1034 136 -974
rect 170 -1034 194 -974
rect 112 -1063 194 -1034
<< nsubdiff >>
rect -102 139 -20 163
rect -102 79 -77 139
rect -43 79 -20 139
rect -102 55 -20 79
<< psubdiffcont >>
rect 136 -1034 170 -974
<< nsubdiffcont >>
rect -77 79 -43 139
<< poly >>
rect 94 14 212 36
rect 94 6 135 14
rect 119 -20 135 6
rect 169 6 212 14
rect 169 -20 185 6
rect 119 -36 185 -20
rect 138 -75 168 -36
rect -80 -349 -50 -188
rect 356 -349 386 -162
rect -80 -365 0 -349
rect -80 -399 -64 -365
rect -30 -399 0 -365
rect -80 -415 0 -399
rect 306 -365 386 -349
rect 306 -399 336 -365
rect 370 -399 386 -365
rect 306 -415 386 -399
rect -80 -774 -50 -696
rect 8 -708 38 -696
rect 8 -724 88 -708
rect 8 -758 38 -724
rect 72 -758 88 -724
rect 8 -774 88 -758
rect 268 -775 298 -696
rect 356 -708 386 -696
rect 356 -724 436 -708
rect 356 -758 386 -724
rect 420 -758 436 -724
rect 356 -774 436 -758
rect -80 -973 -50 -910
rect -96 -989 -30 -973
rect -96 -1023 -80 -989
rect -46 -1023 -30 -989
rect -96 -1039 -30 -1023
rect 268 -1047 298 -910
rect 356 -989 386 -910
rect 356 -1019 416 -989
rect 252 -1063 318 -1047
rect 252 -1097 268 -1063
rect 302 -1097 318 -1063
rect 252 -1113 318 -1097
rect 386 -1168 416 -1019
rect 298 -1707 328 -1652
rect 280 -1723 346 -1707
rect 280 -1757 296 -1723
rect 330 -1757 346 -1723
rect 280 -1773 346 -1757
rect 120 -1793 186 -1777
rect 120 -1827 136 -1793
rect 170 -1827 186 -1793
rect 120 -1833 186 -1827
rect 20 -1863 286 -1833
rect 20 -1905 50 -1863
rect 256 -1905 286 -1863
<< polycont >>
rect 135 -20 169 14
rect -64 -399 -30 -365
rect 336 -399 370 -365
rect 38 -758 72 -724
rect 386 -758 420 -724
rect -80 -1023 -46 -989
rect 268 -1097 302 -1063
rect 296 -1757 330 -1723
rect 136 -1827 170 -1793
<< locali >>
rect -77 300 170 334
rect -77 155 -43 300
rect 136 266 170 300
rect -91 139 -29 155
rect -91 79 -77 139
rect -43 79 -29 139
rect -91 63 -29 79
rect 48 -92 82 58
rect 119 -20 135 14
rect 169 -20 185 14
rect 224 -92 258 58
rect 48 -126 126 -92
rect 180 -126 258 -92
rect -38 -271 -4 -166
rect 310 -271 344 -166
rect -38 -305 92 -271
rect 180 -305 344 -271
rect -80 -399 -64 -365
rect -30 -399 336 -365
rect 370 -399 433 -365
rect -4 -477 84 -443
rect 50 -582 84 -477
rect 398 -582 433 -399
rect -126 -724 -92 -674
rect 222 -724 256 -674
rect -126 -758 38 -724
rect 72 -758 88 -724
rect 222 -758 386 -724
rect 420 -758 436 -724
rect -126 -796 -92 -758
rect 222 -796 256 -758
rect 310 -924 344 -871
rect 120 -958 345 -924
rect 120 -974 186 -958
rect -96 -1023 -80 -989
rect -46 -1023 -30 -989
rect 120 -1034 136 -974
rect 170 -1034 186 -974
rect 120 -1050 186 -1034
rect 120 -1190 157 -1050
rect 252 -1097 268 -1063
rect 302 -1097 318 -1063
rect -77 -1793 -43 -1630
rect 280 -1757 296 -1723
rect 330 -1757 346 -1723
rect -77 -1827 136 -1793
rect 170 -1827 186 -1793
<< viali >>
rect 135 -20 169 14
rect -38 -477 -4 -443
rect -80 -1023 -46 -989
rect 268 -1097 302 -1063
rect 296 -1757 330 -1723
<< metal1 >>
rect -199 308 521 342
rect -171 228 -161 280
rect -109 262 -99 280
rect 136 262 170 308
rect 218 262 268 280
rect -109 228 82 262
rect 258 228 268 262
rect 320 228 330 280
rect 381 75 415 308
rect -57 -26 -47 26
rect 5 20 15 26
rect 343 23 353 75
rect 405 23 415 75
rect 5 14 181 20
rect 5 -20 135 14
rect 169 -20 185 14
rect 5 -26 181 -20
rect -145 -214 -135 -162
rect -83 -214 -73 -162
rect 379 -214 389 -162
rect 441 -214 451 -162
rect 43 -301 53 -249
rect 105 -301 115 -238
rect 191 -301 201 -249
rect 253 -301 263 -249
rect -57 -486 -47 -434
rect 5 -486 15 -434
rect 291 -514 301 -496
rect -199 -548 301 -514
rect 353 -514 363 -496
rect 353 -548 521 -514
rect -38 -586 -4 -548
rect 50 -800 84 -670
rect 136 -722 170 -548
rect 310 -586 344 -548
rect 117 -774 127 -722
rect 179 -774 189 -722
rect 398 -800 432 -670
rect -38 -921 -4 -872
rect 310 -921 344 -872
rect -198 -955 522 -921
rect -92 -989 -34 -983
rect -198 -1023 -80 -989
rect -46 -1023 522 -989
rect -92 -1029 -34 -1023
rect 317 -1057 327 -1051
rect 256 -1063 327 -1057
rect 256 -1097 268 -1063
rect 302 -1097 327 -1063
rect 256 -1103 327 -1097
rect 379 -1103 389 -1051
rect -198 -1165 -125 -1131
rect 510 -1165 522 -1131
rect 117 -1655 127 -1603
rect 179 -1655 189 -1603
rect -198 -1689 -125 -1655
rect 510 -1689 522 -1655
rect 284 -1723 342 -1717
rect -198 -1757 296 -1723
rect 330 -1757 522 -1723
rect 284 -1763 342 -1757
rect 117 -1837 127 -1785
rect 179 -1793 189 -1785
rect 179 -1827 389 -1793
rect 179 -1837 189 -1827
rect 317 -1879 327 -1827
rect 379 -1879 389 -1827
rect 43 -1931 53 -1879
rect 105 -1931 115 -1879
rect 191 -1931 201 -1879
rect 253 -1931 263 -1879
rect -45 -2183 -35 -2131
rect 17 -2183 27 -2131
rect 279 -2183 289 -2131
rect 341 -2183 351 -2131
<< via1 >>
rect -161 228 -109 280
rect 268 228 320 280
rect -47 -26 5 26
rect 353 23 405 75
rect -135 -214 -83 -162
rect 389 -214 441 -162
rect 53 -301 105 -249
rect 201 -301 253 -249
rect -47 -443 5 -434
rect -47 -477 -38 -443
rect -38 -477 -4 -443
rect -4 -477 5 -443
rect -47 -486 5 -477
rect 301 -548 353 -496
rect 127 -774 179 -722
rect 327 -1103 379 -1051
rect 127 -1655 179 -1603
rect 127 -1837 179 -1785
rect 327 -1879 379 -1827
rect 53 -1931 105 -1879
rect 201 -1931 253 -1879
rect -35 -2183 17 -2131
rect 289 -2183 341 -2131
<< metal2 >>
rect -161 280 -109 376
rect -161 218 -109 228
rect 268 280 320 290
rect 429 280 481 376
rect 320 228 481 280
rect 268 218 320 228
rect 301 75 405 85
rect -47 26 5 36
rect -135 -162 -83 -152
rect -135 -985 -83 -214
rect -47 -434 5 -26
rect 301 23 353 75
rect 301 13 405 23
rect -47 -496 5 -486
rect 53 -249 105 -239
rect 53 -632 105 -301
rect -187 -1013 -83 -985
rect 8 -684 105 -632
rect 201 -249 253 -239
rect 201 -632 253 -301
rect 301 -496 353 13
rect 301 -558 353 -548
rect 389 -162 441 -152
rect 201 -684 298 -632
rect -187 -2248 -135 -1013
rect 8 -1871 60 -684
rect 127 -722 179 -712
rect 127 -1603 179 -774
rect 127 -1665 179 -1655
rect 127 -1785 179 -1775
rect 127 -1843 179 -1837
rect 8 -1879 105 -1871
rect 8 -1931 53 -1879
rect 8 -1939 105 -1931
rect 133 -2053 173 -1843
rect 246 -1871 298 -684
rect 389 -985 441 -214
rect 389 -1013 493 -985
rect 201 -1879 298 -1871
rect 253 -1931 298 -1879
rect 327 -1051 379 -1041
rect 327 -1827 379 -1103
rect 327 -1889 379 -1879
rect 201 -1938 298 -1931
rect 441 -1985 493 -1013
rect -35 -2131 17 -2121
rect -35 -2248 17 -2183
rect 127 -2248 179 -2053
rect 289 -2131 341 -2122
rect 289 -2248 341 -2183
rect 441 -2248 494 -1985
use sky130_fd_pr__pfet_01v8_5SMHNA  m1 ~/Desktop/FabRAM/FE/sram130/dido
timestamp 1702473764
transform -1 0 109 0 1 162
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_523TXA  m4 ~/Desktop/FabRAM/FE/sram130/dido
timestamp 1702478055
transform 1 0 -65 0 1 -112
box -109 -112 109 112
use sky130_fd_pr__pfet_01v8_523TXA  m5
timestamp 1702478055
transform -1 0 371 0 1 -112
box -109 -112 109 112
use sky130_fd_pr__nfet_01v8_L8ATA9  m6 ~/Desktop/FabRAM/FE/sram130/dido
timestamp 1702478055
transform -1 0 35 0 1 -2031
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_L8ATA9  m7
timestamp 1702478055
transform 1 0 271 0 1 -2031
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_A6LSUL  m8 ~/Desktop/FabRAM/FE/sram130/common
timestamp 1702483205
transform -1 0 -65 0 1 -842
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m9 ~/Desktop/FabRAM/FE/sram130/common
timestamp 1702483205
transform -1 0 -65 0 1 -628
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m10
timestamp 1702483205
transform 1 0 23 0 1 -628
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_A6LSUL  m11
timestamp 1702483205
transform 1 0 23 0 1 -842
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_A6LSUL  m12
timestamp 1702483205
transform -1 0 283 0 1 -842
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m13
timestamp 1702483205
transform -1 0 283 0 1 -628
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m14
timestamp 1702483205
transform 1 0 371 0 1 -628
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_A6LSUL  m15
timestamp 1702483205
transform 1 0 371 0 1 -842
box -73 -68 73 68
use nand2  nand2_0 ~/Desktop/FabRAM/FE/sram130/nand2
timestamp 1702521001
transform -1 0 510 0 -1 -1040
box 0 91 306 649
use not  not_0 ~/Desktop/FabRAM/FE/sram130/not
timestamp 1702483205
transform -1 0 205 0 -1 -1040
box 0 91 330 649
use sky130_fd_pr__pfet_01v8_5SMHNA  sky130_fd_pr__pfet_01v8_5SMHNA_0
timestamp 1702473764
transform 1 0 197 0 1 162
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_5SMHNA  sky130_fd_pr__pfet_01v8_5SMHNA_1
timestamp 1702473764
transform 1 0 153 0 1 -201
box -109 -162 109 162
<< labels >>
rlabel metal2 -161 324 -109 376 0 BL
rlabel metal2 429 324 481 376 0 BL_
rlabel metal2 -187 -2248 -135 -2196 0 DR
rlabel metal2 -35 -2248 17 -2196 0 DW
rlabel metal2 127 -2248 179 -2196 0 SEL
rlabel metal2 289 -2248 341 -2196 0 DW_
rlabel metal2 441 -2248 493 -2196 0 DR_
rlabel metal1 -199 -548 -165 -514 0 VDD
rlabel metal1 -198 -955 -164 -921 0 VSS
rlabel metal1 -198 -1023 -164 -989 0 PCHG
rlabel metal1 -198 -1165 -164 -1131 0 VSS
rlabel metal1 -198 -1689 -164 -1655 0 VDD
rlabel metal1 -198 -1757 -164 -1723 0 WREN
<< end >>
