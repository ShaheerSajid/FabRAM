magic
tech sky130A
magscale 1 2
timestamp 1702827860
<< nwell >>
rect 0 -236 330 -28
rect 0 -968 328 -760
rect 658 -968 798 -760
rect 1104 -968 1376 -760
rect 1682 -887 1781 -760
rect 1638 -968 1781 -887
rect 2065 -968 2208 -760
rect 2932 -968 3083 -760
rect 1420 -973 1638 -968
<< ndiff >>
rect 3148 -476 3206 -464
rect 3148 -612 3160 -476
rect 3194 -612 3206 -476
rect 3148 -624 3206 -612
<< pdiff >>
rect 3148 -102 3206 -90
rect 3148 -238 3160 -102
rect 3194 -238 3206 -102
rect 3148 -250 3206 -238
<< ndiffc >>
rect 3160 -612 3194 -476
<< pdiffc >>
rect 3160 -238 3194 -102
<< poly >>
rect 206 -92 236 37
rect 2884 -9 2950 7
rect 2884 -43 2900 -9
rect 2934 -43 2950 -9
rect 2884 -59 2950 -43
rect 2900 -64 2930 -59
rect 188 -108 254 -92
rect 188 -142 204 -108
rect 238 -142 254 -108
rect 188 -158 254 -142
rect 3118 -342 3148 -276
rect 3336 -342 3366 -250
rect 2850 -358 2930 -342
rect 2850 -392 2866 -358
rect 2900 -392 2930 -358
rect 2850 -408 2930 -392
rect 3057 -358 3148 -342
rect 3057 -392 3073 -358
rect 3107 -392 3148 -358
rect 3057 -408 3148 -392
rect 3275 -358 3366 -342
rect 3275 -392 3291 -358
rect 3325 -392 3366 -358
rect 3520 -324 3586 -308
rect 3520 -358 3536 -324
rect 3570 -358 3586 -324
rect 3520 -374 3586 -358
rect 3275 -408 3366 -392
rect 2900 -438 2930 -408
rect 3118 -438 3148 -408
rect 3336 -464 3366 -408
rect 3547 -438 3577 -374
rect 1470 -933 1500 -932
rect 1558 -933 1588 -932
rect 1470 -953 1588 -933
rect 1470 -963 1512 -953
rect 1496 -987 1512 -963
rect 1546 -963 1588 -953
rect 1546 -987 1562 -963
rect 1496 -1005 1562 -987
rect 1514 -1009 1544 -1005
<< polycont >>
rect 2900 -43 2934 -9
rect 204 -142 238 -108
rect 2866 -392 2900 -358
rect 3073 -392 3107 -358
rect 3291 -392 3325 -358
rect 3536 -358 3570 -324
rect 1512 -987 1546 -953
<< locali >>
rect 3054 -9 3088 60
rect 2884 -43 2900 -9
rect 2934 -43 3570 -9
rect 3160 -102 3194 -86
rect 188 -142 204 -108
rect 238 -142 436 -108
rect 402 -264 436 -142
rect 2866 -358 2900 -342
rect 2866 -408 2900 -392
rect 2942 -358 2976 -254
rect 3160 -358 3194 -238
rect 2942 -392 3073 -358
rect 3107 -392 3123 -358
rect 3160 -392 3291 -358
rect 3325 -392 3341 -358
rect 2942 -460 2976 -392
rect 3160 -476 3194 -392
rect 3378 -430 3412 -254
rect 3536 -324 3570 -43
rect 3536 -374 3570 -358
rect 3378 -460 3535 -430
rect 3412 -464 3535 -460
rect 1424 -834 1458 -704
rect 1600 -822 1634 -703
rect 3160 -716 3194 -612
rect 3049 -750 3194 -716
rect 1424 -1026 1458 -895
rect 1496 -987 1512 -953
rect 1546 -987 1562 -953
rect 1600 -1026 1634 -910
rect 3049 -954 3083 -750
rect 3049 -988 3128 -954
rect 1424 -1027 1468 -1026
rect 1590 -1027 1634 -1026
rect 1424 -1047 1502 -1027
rect 1556 -1047 1634 -1027
rect 1424 -1061 1468 -1047
rect 1590 -1061 1634 -1047
rect 2558 -1133 2645 -1099
<< viali >>
rect 3160 -238 3194 -102
rect 2866 -392 2900 -358
rect 3160 -612 3194 -476
rect 1424 -704 1458 -670
rect 1600 -703 1634 -669
rect 1512 -987 1546 -953
rect 2645 -1133 2679 -1099
<< metal1 >>
rect 2467 1107 2477 1159
rect 2529 1107 2539 1159
rect 2487 693 2521 1107
rect 2467 641 2477 693
rect 2530 641 2540 693
rect 2854 -28 3024 -27
rect 0 -63 330 -28
rect 2806 -62 3461 -28
rect 2854 -90 2888 -62
rect 3072 -90 3106 -62
rect 3154 -102 3200 -90
rect 3154 -238 3160 -102
rect 3194 -238 3200 -102
rect 3290 -166 3324 -62
rect 3763 -94 3773 -40
rect 3825 -59 3835 -40
rect 3825 -93 4029 -59
rect 3825 -94 3835 -93
rect 3154 -250 3200 -238
rect 0 -283 145 -280
rect 0 -314 83 -283
rect 73 -335 83 -314
rect 135 -335 145 -283
rect 2806 -314 2900 -280
rect 2866 -352 2900 -314
rect 2854 -358 2912 -352
rect 2854 -392 2866 -358
rect 2900 -392 3623 -358
rect 2854 -398 2912 -392
rect 3589 -464 3623 -392
rect 3154 -476 3200 -464
rect 0 -586 330 -552
rect 2806 -586 2854 -552
rect 3154 -612 3160 -476
rect 3194 -612 3200 -476
rect 3154 -624 3200 -612
rect 1405 -704 1415 -652
rect 1467 -704 1477 -652
rect 1405 -710 1477 -704
rect 1580 -703 1590 -651
rect 1642 -703 1652 -651
rect 2854 -653 2888 -624
rect 3072 -653 3106 -624
rect 3290 -653 3324 -548
rect 2854 -687 3325 -653
rect 1580 -709 1652 -703
rect 0 -794 328 -760
rect 658 -794 798 -760
rect 1104 -794 1424 -760
rect 1458 -794 1735 -760
rect 2065 -794 2208 -760
rect 2932 -794 3083 -760
rect 772 -988 806 -794
rect 3878 -827 4028 -793
rect 1677 -947 1687 -922
rect 1500 -953 1687 -947
rect 1070 -987 1512 -953
rect 1546 -974 1687 -953
rect 1739 -974 1749 -922
rect 2146 -968 2156 -916
rect 2208 -968 2218 -916
rect 3719 -968 3736 -916
rect 3788 -968 3798 -916
rect 1546 -981 1749 -974
rect 1546 -987 1558 -981
rect 318 -1012 328 -1002
rect 0 -1046 328 -1012
rect 318 -1054 328 -1046
rect 380 -1054 390 -1002
rect 658 -1046 738 -1012
rect 1070 -1046 1104 -987
rect 1500 -993 1558 -987
rect 1707 -1034 1735 -1012
rect 704 -1099 738 -1046
rect 1596 -1068 1735 -1034
rect 2029 -1058 2208 -1024
rect 2932 -1047 2997 -1012
rect 3719 -1046 3753 -968
rect 3878 -1003 3912 -827
rect 704 -1133 798 -1099
rect 2146 -1148 2156 -1096
rect 2208 -1148 2218 -1096
rect 2633 -1099 2691 -1093
rect 2963 -1099 2997 -1047
rect 3857 -1055 3867 -1003
rect 3919 -1055 3929 -1003
rect 2633 -1133 2645 -1099
rect 2679 -1133 3083 -1099
rect 2633 -1139 2691 -1133
rect 2963 -1192 2997 -1133
rect 2963 -1245 2973 -1192
rect 3025 -1245 3035 -1192
rect 0 -1318 328 -1284
rect 658 -1318 798 -1284
rect 1104 -1318 1735 -1284
rect 2065 -1318 2208 -1284
rect 2932 -1318 3083 -1284
<< via1 >>
rect 2477 1107 2529 1159
rect 2477 641 2530 693
rect 3773 -94 3825 -40
rect 83 -335 135 -283
rect 1415 -670 1467 -652
rect 1415 -704 1424 -670
rect 1424 -704 1458 -670
rect 1458 -704 1467 -670
rect 1590 -669 1642 -651
rect 1590 -703 1600 -669
rect 1600 -703 1634 -669
rect 1634 -703 1642 -669
rect 1687 -974 1739 -922
rect 2156 -968 2208 -916
rect 3736 -968 3788 -916
rect 328 -1054 380 -1002
rect 2156 -1148 2208 -1096
rect 3867 -1055 3919 -1003
rect 2973 -1245 3025 -1192
<< metal2 >>
rect 2477 1159 2529 1306
rect 2477 1097 2529 1107
rect 3346 979 3398 1306
rect 1424 945 3398 979
rect 83 -283 135 -273
rect 83 -345 135 -335
rect 93 -1105 127 -345
rect 1424 -642 1458 945
rect 3936 870 3988 1306
rect 1600 836 3988 870
rect 1600 -641 1634 836
rect 2477 693 2530 703
rect 2530 641 3912 665
rect 2477 631 3912 641
rect 3773 -40 3825 -30
rect 3773 -104 3825 -94
rect 1415 -652 1467 -642
rect 1415 -714 1467 -704
rect 1590 -651 1642 -641
rect 1590 -713 1642 -703
rect 3782 -811 3816 -104
rect 1739 -845 3816 -811
rect 1739 -912 1773 -845
rect 3878 -906 3912 631
rect 1687 -922 1773 -912
rect 1739 -974 1773 -922
rect 1687 -984 1773 -974
rect 2156 -916 2208 -906
rect 3736 -916 3912 -906
rect 2208 -968 3736 -934
rect 3788 -940 3912 -916
rect 2156 -978 2208 -968
rect 3736 -978 3788 -968
rect 328 -1002 380 -992
rect 3867 -1003 3919 -993
rect 380 -1046 3867 -1012
rect 328 -1064 380 -1054
rect 3867 -1065 3919 -1055
rect 2156 -1096 2208 -1086
rect 93 -1139 2156 -1105
rect 2156 -1158 2208 -1148
rect 2973 -1192 3025 -1182
rect 2973 -1318 3025 -1245
use del_cell  del_cell_0
timestamp 1702826916
transform 1 0 496 0 1 1
box -166 -1 2310 557
use del_cell  del_cell_1
timestamp 1702826916
transform 1 0 496 0 1 -585
box -166 -1 2310 557
use sky130_fd_pr__nfet_01v8_BBXUYH  m1
timestamp 1702809544
transform 1 0 2915 0 1 -544
box -73 -106 73 106
use sky130_fd_pr__pfet_01v8_5C6TXA  m2
timestamp 1702809544
transform 1 0 2915 0 1 -170
box -109 -142 109 142
use sky130_fd_pr__pfet_01v8_5C6TXA  m3
timestamp 1702809544
transform 1 0 3133 0 1 -170
box -109 -142 109 142
use sky130_fd_pr__nfet_01v8_BBXUYH  m4
timestamp 1702809544
transform 1 0 3133 0 1 -544
box -73 -106 73 106
use sky130_fd_pr__pfet_01v8_4Y88KP  m5
timestamp 1702809649
transform 1 0 3351 0 1 -208
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_A6LSUL  m6
timestamp 1702809544
transform 1 0 3351 0 1 -506
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_BBXUYH  m7
timestamp 1702809544
transform 1 0 3562 0 1 -544
box -73 -106 73 106
use sky130_fd_pr__pfet_01v8_4Y88KP  m8
timestamp 1702809649
transform -1 0 1485 0 1 -864
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m9
timestamp 1702809649
transform 1 0 1573 0 1 -864
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m10
timestamp 1702809649
transform 1 0 1529 0 1 -1077
box -109 -104 109 104
use nand2_f  nand2_f_0 ~/Desktop/FabRAM/FE/sram130/nand2
timestamp 1702826916
transform 1 0 3083 0 1 -1456
box 0 138 306 696
use nand2_f  nand2_f_1
timestamp 1702826916
transform 1 0 798 0 1 -1456
box 0 138 306 696
use nand3_f  nand3_f_0 ~/Desktop/FabRAM/FE/sram130/nand3
timestamp 1702826916
transform 1 0 2208 0 1 -1456
box 0 138 394 696
use not_f  not_f_0 ~/Desktop/FabRAM/FE/sram130/not
timestamp 1702826916
transform 1 0 0 0 1 -138
box 0 138 330 696
use not_f  not_f_1
timestamp 1702826916
transform 1 0 2806 0 1 -137
box 0 138 330 696
use not_f  not_f_2
timestamp 1702826916
transform 1 0 3389 0 1 -1456
box 0 138 330 696
use not_f  not_f_3
timestamp 1702826916
transform 1 0 328 0 1 -1456
box 0 138 330 696
use not_f  not_f_4
timestamp 1702826916
transform 1 0 1735 0 1 -1456
box 0 138 330 696
use not_f  not_f_5
timestamp 1702826916
transform 1 0 2602 0 1 -1456
box 0 138 330 696
<< end >>
