.title sram_gen
.subckt bit_cell VDD VSS WL BL BL_
X0 Q Q_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X1 Q_ Q VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X2 Q Q_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 Q_ Q VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 Q WL BL VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
X5 Q_ WL BL_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
.ends bit_cell

.subckt dmy_cell VDD VSS WL BL BL_
X0 Q VSS VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X1 Q_ VDD VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X2 Q VSS VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 Q_ VDD VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 Q WL BL VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
X5 Q_ WL BL_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
.ends dmy_cell

.subckt in_reg VDD VSS clk D Q
X0 net3 clk VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X8 net3 clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 net4 net2 net5 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X10 Din net2 net1 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 net55 Q VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X13 net55 Q VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 net2 net3 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X11 net2 net3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X5 Din net3 net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X15 net4 net3 net5 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 Q net5 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X9 Q net5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X6 net11 net4 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X12 net11 net4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X7 net4 net1 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X14 net4 net1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X16 net11 net2 net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X17 net11 net3 net1 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X18 net55 net3 net5 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X19 net55 net2 net5 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X20 D_ D VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X21 D_ D VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X22 Din D_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X23 Din D_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
.ends in_reg

.subckt se_cell VDD VSS SAEN BL BL_ SB
X0 net1 SAEN VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.84
X1 diff1 BL_ net1 net1 sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X2 diff2 BL net1 net1 sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X3 diff1 diff1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 diff2 diff1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X5 diff2_ diff2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X6 diff2_ diff2 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=2
X7 SB_ diff2_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X8 SB_ diff2_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=2
X9 SB_w Q_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X10 Q_ SB_w VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X11 SB_w Q_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X12 Q_ SB_w VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X13 SB_w SAEN SB_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
X14 Q_ SAEN diff2_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
X15 SB SB_w VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X16 SB SB_w VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
.ends se_cell

.subckt not VDD VSS A B
X0 B A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 B A VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends not

.subckt notdel VDD VSS A B
X0 B A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.84
X1 B A VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends notdel

.subckt nand2 VDD VSS A B Y
X0 Y A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 Y B VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 Y B net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X3 net1 A VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends nand2

.subckt nand3 VDD VSS A B C Y
X0 Y A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 Y B VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 Y C VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 Y A net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X4 net1 B net2 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X5 net2 C VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends nand3

.subckt nand4 VDD VSS A B C D Y
X0 Y A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 Y B VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 Y C VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 Y D VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 Y D net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X5 net1 B net2 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X6 net2 C net3 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X7 net3 A VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends nand4

.subckt dec_2to4 VDD VSS A1 A0 Y0 Y1 Y2 Y3
X0 VDD VSS A1 A_1 not
X1 VDD VSS A0 A_0 not
X2 VDD VSS A_1 A_0 Y0_ nand2
X3 VDD VSS A_1 A0 Y1_ nand2
X4 VDD VSS A1 A_0 Y2_ nand2
X5 VDD VSS A1 A0 Y3_ nand2
X6 VDD VSS Y0_ Y0 not
X7 VDD VSS Y1_ Y1 not
X8 VDD VSS Y2_ Y2 not
X9 VDD VSS Y3_ Y3 not
.ends dec_2to4

.subckt dec_3to6 VDD VSS A2 A1 A0 Y0 Y1 Y2 Y3 Y4 Y5
X0 VDD VSS A2 Y4 not
X1 VDD VSS Y4 Y5 not
X2 VDD VSS A1 A0 Y0 Y1 Y2 Y3 dec_2to4
.ends dec_3to6

.subckt row_dec32 VDD VSS A0 A1 A2 A3 A4 DC0 DC1 DC2 DC3 DC4 DC5 DC6 DC7 DC8 DC9 DC10 DC11 DC12 DC13 DC14 DC15 DC16 DC17 DC18 DC19 DC20 DC21 DC22 DC23 DC24 DC25 DC26 DC27 DC28 DC29 DC30 DC31
X0 VDD VSS A1 A0 Y0 Y1 Y2 Y3 dec_2to4
X1 VDD VSS A4 A3 A2 Y4 Y5 Y6 Y7 Y8 Y9 dec_3to6
X2 VDD VSS Y0 Y4 Y8 DC_0 nand3
X3 VDD VSS Y1 Y4 Y8 DC_1 nand3
X4 VDD VSS Y2 Y4 Y8 DC_2 nand3
X5 VDD VSS Y3 Y4 Y8 DC_3 nand3
X6 VDD VSS Y0 Y5 Y8 DC_4 nand3
X7 VDD VSS Y1 Y5 Y8 DC_5 nand3
X8 VDD VSS Y2 Y5 Y8 DC_6 nand3
X9 VDD VSS Y3 Y5 Y8 DC_7 nand3
X10 VDD VSS Y0 Y6 Y8 DC_8 nand3
X11 VDD VSS Y1 Y6 Y8 DC_9 nand3
X12 VDD VSS Y2 Y6 Y8 DC_10 nand3
X13 VDD VSS Y3 Y6 Y8 DC_11 nand3
X14 VDD VSS Y0 Y7 Y8 DC_12 nand3
X15 VDD VSS Y1 Y7 Y8 DC_13 nand3
X16 VDD VSS Y2 Y7 Y8 DC_14 nand3
X17 VDD VSS Y3 Y7 Y8 DC_15 nand3
X18 VDD VSS Y0 Y4 Y9 DC_16 nand3
X19 VDD VSS Y1 Y4 Y9 DC_17 nand3
X20 VDD VSS Y2 Y4 Y9 DC_18 nand3
X21 VDD VSS Y3 Y4 Y9 DC_19 nand3
X22 VDD VSS Y0 Y5 Y9 DC_20 nand3
X23 VDD VSS Y1 Y5 Y9 DC_21 nand3
X24 VDD VSS Y2 Y5 Y9 DC_22 nand3
X25 VDD VSS Y3 Y5 Y9 DC_23 nand3
X26 VDD VSS Y0 Y6 Y9 DC_24 nand3
X27 VDD VSS Y1 Y6 Y9 DC_25 nand3
X28 VDD VSS Y2 Y6 Y9 DC_26 nand3
X29 VDD VSS Y3 Y6 Y9 DC_27 nand3
X30 VDD VSS Y0 Y7 Y9 DC_28 nand3
X31 VDD VSS Y1 Y7 Y9 DC_29 nand3
X32 VDD VSS Y2 Y7 Y9 DC_30 nand3
X33 VDD VSS Y3 Y7 Y9 DC_31 nand3
X34 VDD VSS DC_0 DC0 not
X35 VDD VSS DC_1 DC1 not
X36 VDD VSS DC_2 DC2 not
X37 VDD VSS DC_3 DC3 not
X38 VDD VSS DC_4 DC4 not
X39 VDD VSS DC_5 DC5 not
X40 VDD VSS DC_6 DC6 not
X41 VDD VSS DC_7 DC7 not
X42 VDD VSS DC_8 DC8 not
X43 VDD VSS DC_9 DC9 not
X44 VDD VSS DC_10 DC10 not
X45 VDD VSS DC_11 DC11 not
X46 VDD VSS DC_12 DC12 not
X47 VDD VSS DC_13 DC13 not
X48 VDD VSS DC_14 DC14 not
X49 VDD VSS DC_15 DC15 not
X50 VDD VSS DC_16 DC16 not
X51 VDD VSS DC_17 DC17 not
X52 VDD VSS DC_18 DC18 not
X53 VDD VSS DC_19 DC19 not
X54 VDD VSS DC_20 DC20 not
X55 VDD VSS DC_21 DC21 not
X56 VDD VSS DC_22 DC22 not
X57 VDD VSS DC_23 DC23 not
X58 VDD VSS DC_24 DC24 not
X59 VDD VSS DC_25 DC25 not
X60 VDD VSS DC_26 DC26 not
X61 VDD VSS DC_27 DC27 not
X62 VDD VSS DC_28 DC28 not
X63 VDD VSS DC_29 DC29 not
X64 VDD VSS DC_30 DC30 not
X65 VDD VSS DC_31 DC31 not
.ends row_dec32

.subckt row_driver VDD VSS WLEN A B
X0 VDD VSS A WLEN net1 nand2
X1 B net1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X2 B net1 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
.ends row_driver

.subckt rd_arr_32 VDD VSS WLEN DC0 DC1 DC2 DC3 DC4 DC5 DC6 DC7 DC8 DC9 DC10 DC11 DC12 DC13 DC14 DC15 DC16 DC17 DC18 DC19 DC20 DC21 DC22 DC23 DC24 DC25 DC26 DC27 DC28 DC29 DC30 DC31 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31
X0 VDD VSS WLEN DC0 WL0 row_driver
X1 VDD VSS WLEN DC1 WL1 row_driver
X2 VDD VSS WLEN DC2 WL2 row_driver
X3 VDD VSS WLEN DC3 WL3 row_driver
X4 VDD VSS WLEN DC4 WL4 row_driver
X5 VDD VSS WLEN DC5 WL5 row_driver
X6 VDD VSS WLEN DC6 WL6 row_driver
X7 VDD VSS WLEN DC7 WL7 row_driver
X8 VDD VSS WLEN DC8 WL8 row_driver
X9 VDD VSS WLEN DC9 WL9 row_driver
X10 VDD VSS WLEN DC10 WL10 row_driver
X11 VDD VSS WLEN DC11 WL11 row_driver
X12 VDD VSS WLEN DC12 WL12 row_driver
X13 VDD VSS WLEN DC13 WL13 row_driver
X14 VDD VSS WLEN DC14 WL14 row_driver
X15 VDD VSS WLEN DC15 WL15 row_driver
X16 VDD VSS WLEN DC16 WL16 row_driver
X17 VDD VSS WLEN DC17 WL17 row_driver
X18 VDD VSS WLEN DC18 WL18 row_driver
X19 VDD VSS WLEN DC19 WL19 row_driver
X20 VDD VSS WLEN DC20 WL20 row_driver
X21 VDD VSS WLEN DC21 WL21 row_driver
X22 VDD VSS WLEN DC22 WL22 row_driver
X23 VDD VSS WLEN DC23 WL23 row_driver
X24 VDD VSS WLEN DC24 WL24 row_driver
X25 VDD VSS WLEN DC25 WL25 row_driver
X26 VDD VSS WLEN DC26 WL26 row_driver
X27 VDD VSS WLEN DC27 WL27 row_driver
X28 VDD VSS WLEN DC28 WL28 row_driver
X29 VDD VSS WLEN DC29 WL29 row_driver
X30 VDD VSS WLEN DC30 WL30 row_driver
X31 VDD VSS WLEN DC31 WL31 row_driver
.ends rd_arr_32

.subckt col_dec1 VDD VSS DC0
X0 DC0 VDD VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X1 DC0 VDD VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
.ends col_dec1

.subckt dido VDD VSS PCHG WREN SEL BL BL_ DW DW_ DR DR_
X0 BL_ net6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 BL net6 BL_ VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 BL net6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 net6 net5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 net6 net5 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X5 net5 PCHG VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X6 net5 PCHG VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X7 BL_ net3 DR_ VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X8 DR net3 BL VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X9 net4 SEL VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X10 BL net2 DW VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X11 DW_ net2 BL_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X12 net4 SEL VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X13 net3 net4 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X14 net3 net4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X15 VDD VSS net4 WREN net1 nand2
X16 VDD VSS net1 net2 not
.ends dido

.subckt dido_arr_4 VDD VSS PCHG WREN SEL0 SEL1 SEL2 SEL3 BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 DW0 DW_0 DW1 DW_1 DW2 DW_2 DW3 DW_3 DR0 DR_0 DR1 DR_1 DR2 DR_2 DR3 DR_3
X0 VDD VSS PCHG WREN SEL0 BL0 BL_0 DW0 DW_0 DR0 DR_0 dido
X1 VDD VSS PCHG WREN SEL1 BL1 BL_1 DW1 DW_1 DR1 DR_1 dido
X2 VDD VSS PCHG WREN SEL2 BL2 BL_2 DW2 DW_2 DR2 DR_2 dido
X3 VDD VSS PCHG WREN SEL3 BL3 BL_3 DW3 DW_3 DR3 DR_3 dido
.ends dido_arr_4

.subckt write_driver VDD VSS WREN Din DW DW_
X0 en_ WREN VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 en_ WREN VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X4 d_ Din VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X5 d_ Din VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X6 net1 Din VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X7 DW_ en_ net1 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X8 DW_ WREN net2 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
X9 net2 Din VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
X10 net3 d_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X11 DW en_ net3 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X12 DW WREN net4 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
X13 net4 d_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
.ends write_driver

.subckt del10 VDD VSS A B
X0 VDD VSS A net1 notdel
X1 VDD VSS net1 net2 notdel
X2 VDD VSS net2 net3 notdel
X3 VDD VSS net3 net4 notdel
X4 VDD VSS net4 net5 notdel
X5 VDD VSS net5 net6 notdel
X6 VDD VSS net6 net7 notdel
X7 VDD VSS net7 net8 notdel
X8 VDD VSS net8 net9 notdel
X9 VDD VSS net9 net10 notdel
X10 VDD VSS net10 net11 notdel
X11 VDD VSS A net11 net12 nand2
X12 VDD VSS net12 B not
.ends del10

.subckt ctrl VDD VSS clk cs write DBL DBL_ WREN PCHG WLEN SAEN
X0 clk_ clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 clk_ clk VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X2 WLENP clk_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 WLENP clk_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X4 VDD VSS write WREN_ not
X8 PCHG clk_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X9 PCHG clk_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
X10 DBL_ PCHG VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X11 DBL PCHG DBL_ VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X12 DBL PCHG VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X13 VDD VSS cs WLENP WLENPP nand2
X21 WLEN WLENPP VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X22 WLEN WLENPP VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
X15 VDD VSS DBL_ RBL not
X16 VDD VSS WLEN RBL SAEN_ nand2
X17 SAEN SAEN_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X18 SAEN SAEN_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
X19 WREN WREN_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X20 WREN WREN_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
.ends ctrl

.subckt input_reg6 VDD VSS clk D0 D1 D2 D3 D4 D5 Q0 Q1 Q2 Q3 Q4 Q5
X0 VDD VSS clk D0 Q0 in_reg
X1 VDD VSS clk D1 Q1 in_reg
X2 VDD VSS clk D2 Q2 in_reg
X3 VDD VSS clk D3 Q3 in_reg
X4 VDD VSS clk D4 Q4 in_reg
X5 VDD VSS clk D5 Q5 in_reg
.ends input_reg6

.subckt datain_reg4 VDD VSS clk WREN din0 din1 din2 din3 DW0 DW_0 DW1 DW_1 DW2 DW_2 DW3 DW_3
X0 VDD VSS clk din0 din_r0 in_reg
X1 VDD VSS clk din1 din_r1 in_reg
X2 VDD VSS clk din2 din_r2 in_reg
X3 VDD VSS clk din3 din_r3 in_reg
X4 VDD VSS WREN din_r0 DW0 DW_0 write_driver
X8 VDD VSS WREN din_r1 DW1 DW_1 write_driver
X12 VDD VSS WREN din_r2 DW2 DW_2 write_driver
X16 VDD VSS WREN din_r3 DW3 DW_3 write_driver
.ends datain_reg4

.subckt bit_arr_4 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL
X0 VDD VSS WL BL0 BL_0 bit_cell
X1 VDD VSS WL BL1 BL_1 bit_cell
X2 VDD VSS WL BL2 BL_2 bit_cell
X3 VDD VSS WL BL3 BL_3 bit_cell
.ends bit_arr_4

.subckt dmy_arr_32 VDD VSS WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 DBL DBL_
X0 VDD VSS WL0 DBL DBL_ dmy_cell
X1 VDD VSS WL1 DBL DBL_ dmy_cell
X2 VDD VSS WL2 DBL DBL_ dmy_cell
X3 VDD VSS WL3 DBL DBL_ dmy_cell
X4 VDD VSS WL4 DBL DBL_ dmy_cell
X5 VDD VSS WL5 DBL DBL_ dmy_cell
X6 VDD VSS WL6 DBL DBL_ dmy_cell
X7 VDD VSS WL7 DBL DBL_ dmy_cell
X8 VDD VSS WL8 DBL DBL_ dmy_cell
X9 VDD VSS WL9 DBL DBL_ dmy_cell
X10 VDD VSS WL10 DBL DBL_ dmy_cell
X11 VDD VSS WL11 DBL DBL_ dmy_cell
X12 VDD VSS WL12 DBL DBL_ dmy_cell
X13 VDD VSS WL13 DBL DBL_ dmy_cell
X14 VDD VSS WL14 DBL DBL_ dmy_cell
X15 VDD VSS WL15 DBL DBL_ dmy_cell
X16 VDD VSS WL16 DBL DBL_ dmy_cell
X17 VDD VSS WL17 DBL DBL_ dmy_cell
X18 VDD VSS WL18 DBL DBL_ dmy_cell
X19 VDD VSS WL19 DBL DBL_ dmy_cell
X20 VDD VSS WL20 DBL DBL_ dmy_cell
X21 VDD VSS WL21 DBL DBL_ dmy_cell
X22 VDD VSS WL22 DBL DBL_ dmy_cell
X23 VDD VSS WL23 DBL DBL_ dmy_cell
X24 VDD VSS WL24 DBL DBL_ dmy_cell
X25 VDD VSS WL25 DBL DBL_ dmy_cell
X26 VDD VSS WL26 DBL DBL_ dmy_cell
X27 VDD VSS WL27 DBL DBL_ dmy_cell
X28 VDD VSS WL28 DBL DBL_ dmy_cell
X29 VDD VSS WL29 DBL DBL_ dmy_cell
X30 VDD VSS WL30 DBL DBL_ dmy_cell
X31 VDD VSS WL31 DBL DBL_ dmy_cell
.ends dmy_arr_32

.subckt se_arr_4 VDD VSS SAEN BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 SB0 SB1 SB2 SB3
X0 VDD VSS SAEN BL0 BL_0 SB0 se_cell
X1 VDD VSS SAEN BL1 BL_1 SB1 se_cell
X2 VDD VSS SAEN BL2 BL_2 SB2 se_cell
X3 VDD VSS SAEN BL3 BL_3 SB3 se_cell
.ends se_arr_4

.subckt mat_arr_4 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31
X0 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL0 bit_arr_4
X1 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL1 bit_arr_4
X2 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL2 bit_arr_4
X3 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL3 bit_arr_4
X4 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL4 bit_arr_4
X5 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL5 bit_arr_4
X6 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL6 bit_arr_4
X7 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL7 bit_arr_4
X8 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL8 bit_arr_4
X9 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL9 bit_arr_4
X10 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL10 bit_arr_4
X11 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL11 bit_arr_4
X12 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL12 bit_arr_4
X13 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL13 bit_arr_4
X14 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL14 bit_arr_4
X15 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL15 bit_arr_4
X16 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL16 bit_arr_4
X17 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL17 bit_arr_4
X18 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL18 bit_arr_4
X19 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL19 bit_arr_4
X20 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL20 bit_arr_4
X21 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL21 bit_arr_4
X22 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL22 bit_arr_4
X23 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL23 bit_arr_4
X24 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL24 bit_arr_4
X25 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL25 bit_arr_4
X26 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL26 bit_arr_4
X27 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL27 bit_arr_4
X28 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL28 bit_arr_4
X29 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL29 bit_arr_4
X30 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL30 bit_arr_4
X31 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL31 bit_arr_4
.ends mat_arr_4

.subckt sram32x4 VDD VSS clk addr0 addr1 addr2 addr3 addr4 din0 din1 din2 din3 Q0 Q1 Q2 Q3 w_en cs
X0 VDD VSS clk addr0 addr1 addr2 addr3 addr4 w_en A0 A1 A2 A3 A4 write input_reg6
X1 VDD VSS A0 A1 A2 A3 A4 DC0 DC1 DC2 DC3 DC4 DC5 DC6 DC7 DC8 DC9 DC10 DC11 DC12 DC13 DC14 DC15 DC16 DC17 DC18 DC19 DC20 DC21 DC22 DC23 DC24 DC25 DC26 DC27 DC28 DC29 DC30 DC31 row_dec32
X2 VDD VSS WLEN DC0 DC1 DC2 DC3 DC4 DC5 DC6 DC7 DC8 DC9 DC10 DC11 DC12 DC13 DC14 DC15 DC16 DC17 DC18 DC19 DC20 DC21 DC22 DC23 DC24 DC25 DC26 DC27 DC28 DC29 DC30 DC31 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 rd_arr_32
X3 VDD VSS SEL0 col_dec1
X4 VDD VSS PCHG WREN SEL0 SEL0 SEL0 SEL0 BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 DW0 DW_0 DW1 DW_1 DW2 DW_2 DW3 DW_3 DR0 DR_0 DR1 DR_1 DR2 DR_2 DR3 DR_3 dido_arr_4
X5 VDD VSS clk WREN din0 din1 din2 din3 DW0 DW_0 DW1 DW_1 DW2 DW_2 DW3 DW_3 datain_reg4
X6 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 mat_arr_4
X7 VDD VSS SAEN DR0 DR_0 DR1 DR_1 DR2 DR_2 DR3 DR_3 Q0 Q1 Q2 Q3 se_arr_4
X8 VDD VSS clk cs write DBL DBL_ WREN PCHG WLEN SAEN ctrl
X9 VDD VSS WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 DBL DBL_ dmy_arr_32
.ends sram32x4

