magic
tech sky130A
magscale 1 2
timestamp 1703660268
<< metal1 >>
rect 2179 -217 2213 0
rect 2179 -251 2300 -217
rect 1163 -586 1173 -564
rect 831 -620 1173 -586
rect 1229 -620 1239 -564
rect 1257 -1282 1267 -1260
rect 831 -1316 1267 -1282
rect 1323 -1316 1333 -1260
<< via1 >>
rect 1173 -620 1229 -564
rect 1267 -1316 1323 -1260
<< metal2 >>
rect 1173 783 1229 793
rect 1173 -564 1229 727
rect 1173 -638 1229 -620
rect 1267 657 1323 667
rect 1267 -1260 1323 601
rect 1267 -1327 1323 -1316
<< via2 >>
rect 1173 727 1229 783
rect 1267 601 1323 657
<< metal3 >>
rect 1163 783 2289 788
rect 1163 727 1173 783
rect 1229 727 2289 783
rect 1163 722 2289 727
rect 1257 657 2289 662
rect 1257 601 1267 657
rect 1323 601 2289 657
rect 1257 596 2289 601
use col_dec2_f  col_dec2_f_0
timestamp 1703656013
transform 1 0 0 0 1 0
box 0 0 2301 1165
<< end >>
