magic
tech sky130A
magscale 1 2
timestamp 1703822710
<< nwell >>
rect 271 350 841 558
<< nmos >>
rect 365 63 395 147
rect 453 63 483 147
rect 541 63 571 147
rect 629 63 659 147
rect 717 63 747 147
<< pmos >>
rect 365 412 395 496
rect 453 412 483 496
rect 541 412 571 496
rect 629 412 659 496
rect 717 412 747 496
<< ndiff >>
rect 307 122 365 147
rect 307 88 319 122
rect 353 88 365 122
rect 307 63 365 88
rect 395 122 453 147
rect 395 88 407 122
rect 441 88 453 122
rect 395 63 453 88
rect 483 122 541 147
rect 483 88 495 122
rect 529 88 541 122
rect 483 63 541 88
rect 571 122 629 147
rect 571 88 583 122
rect 617 88 629 122
rect 571 63 629 88
rect 659 122 717 147
rect 659 88 671 122
rect 705 88 717 122
rect 659 63 717 88
rect 747 122 805 147
rect 747 88 759 122
rect 793 88 805 122
rect 747 63 805 88
<< pdiff >>
rect 307 471 365 496
rect 307 437 319 471
rect 353 437 365 471
rect 307 412 365 437
rect 395 471 453 496
rect 395 437 407 471
rect 441 437 453 471
rect 395 412 453 437
rect 483 471 541 496
rect 483 437 495 471
rect 529 437 541 471
rect 483 412 541 437
rect 571 471 629 496
rect 571 437 583 471
rect 617 437 629 471
rect 571 412 629 437
rect 659 471 717 496
rect 659 437 671 471
rect 705 437 717 471
rect 659 412 717 437
rect 747 471 805 496
rect 747 437 759 471
rect 793 437 805 471
rect 747 412 805 437
<< ndiffc >>
rect 319 88 353 122
rect 407 88 441 122
rect 495 88 529 122
rect 583 88 617 122
rect 671 88 705 122
rect 759 88 793 122
<< pdiffc >>
rect 319 437 353 471
rect 407 437 441 471
rect 495 437 529 471
rect 583 437 617 471
rect 671 437 705 471
rect 759 437 793 471
<< poly >>
rect 365 496 395 522
rect 453 496 483 522
rect 541 496 571 522
rect 629 496 659 522
rect 717 496 747 522
rect 365 324 395 412
rect 312 306 395 324
rect 453 306 483 412
rect 541 306 571 412
rect 629 306 659 412
rect 717 306 747 412
rect 312 272 322 306
rect 356 272 747 306
rect 312 256 395 272
rect 365 147 395 256
rect 453 147 483 272
rect 541 147 571 272
rect 629 147 659 272
rect 717 147 747 272
rect 365 37 395 63
rect 453 37 483 63
rect 541 37 571 63
rect 629 37 659 63
rect 717 37 747 63
<< polycont >>
rect 322 272 356 306
<< locali >>
rect 319 471 353 500
rect 319 408 353 437
rect 407 471 441 500
rect 407 358 441 437
rect 495 471 529 500
rect 495 408 529 437
rect 583 471 617 500
rect 583 358 617 437
rect 671 471 705 500
rect 671 408 705 437
rect 759 471 793 500
rect 759 358 793 437
rect 407 323 793 358
rect 759 306 793 323
rect 305 272 322 306
rect 356 272 372 306
rect 759 220 793 272
rect 407 185 793 220
rect 319 122 353 151
rect 319 59 353 88
rect 407 122 441 185
rect 407 59 441 88
rect 495 122 529 151
rect 495 59 529 88
rect 583 122 617 185
rect 583 59 617 88
rect 671 122 705 151
rect 671 59 705 88
rect 759 122 793 185
rect 759 59 793 88
<< viali >>
rect 319 437 353 471
rect 407 437 441 471
rect 495 437 529 471
rect 583 437 617 471
rect 671 437 705 471
rect 759 437 793 471
rect 322 272 356 306
rect 759 272 793 306
rect 319 88 353 122
rect 407 88 441 122
rect 495 88 529 122
rect 583 88 617 122
rect 671 88 705 122
rect 759 88 793 122
<< metal1 >>
rect 272 524 841 558
rect 319 496 353 524
rect 495 496 529 524
rect 671 496 705 524
rect 313 471 359 496
rect 313 437 319 471
rect 353 437 359 471
rect 313 412 359 437
rect 401 471 447 496
rect 401 437 407 471
rect 441 437 447 471
rect 401 412 447 437
rect 489 471 535 496
rect 489 437 495 471
rect 529 437 535 471
rect 489 412 535 437
rect 577 471 623 496
rect 577 437 583 471
rect 617 437 623 471
rect 577 412 623 437
rect 665 471 711 496
rect 665 437 671 471
rect 705 437 711 471
rect 665 412 711 437
rect 753 471 799 496
rect 753 437 759 471
rect 793 437 799 471
rect 753 412 799 437
rect 310 306 368 312
rect 0 301 322 306
rect 0 249 10 301
rect 62 272 322 301
rect 356 272 368 306
rect 62 249 72 272
rect 310 266 368 272
rect 747 306 805 312
rect 995 306 1005 328
rect 747 272 759 306
rect 793 272 1005 306
rect 1061 272 1071 328
rect 747 266 805 272
rect 2189 169 2223 665
rect 313 122 359 147
rect 313 88 319 122
rect 353 88 359 122
rect 313 63 359 88
rect 401 122 447 147
rect 401 88 407 122
rect 441 88 447 122
rect 401 63 447 88
rect 489 122 535 147
rect 489 88 495 122
rect 529 88 535 122
rect 489 63 535 88
rect 577 122 623 147
rect 577 88 583 122
rect 617 88 623 122
rect 577 63 623 88
rect 665 122 711 147
rect 665 88 671 122
rect 705 88 711 122
rect 665 63 711 88
rect 753 122 799 147
rect 2189 135 2299 169
rect 753 88 759 122
rect 793 88 799 122
rect 753 63 799 88
rect 319 34 353 63
rect 495 34 529 63
rect 671 34 705 63
rect 272 0 841 34
<< via1 >>
rect 10 249 62 301
rect 1005 272 1061 328
<< metal2 >>
rect 10 301 63 665
rect 62 249 63 301
rect 1005 535 1061 545
rect 1005 328 1061 479
rect 1005 262 1061 272
rect 10 239 62 249
<< via2 >>
rect 1005 479 1061 535
<< metal3 >>
rect 995 535 2299 540
rect 995 479 1005 535
rect 1061 479 2299 535
rect 995 474 2299 479
<< end >>
