magic
tech sky130A
magscale 1 2
timestamp 1703586424
<< nwell >>
rect 0 488 876 696
<< pwell >>
rect 10 175 866 311
<< nmos >>
rect 94 201 124 285
rect 182 201 212 285
rect 400 201 430 285
rect 488 201 518 285
rect 576 201 606 285
rect 664 201 694 285
rect 752 201 782 285
<< pmos >>
rect 94 550 124 634
rect 182 550 212 634
rect 400 550 430 634
rect 488 550 518 634
rect 576 550 606 634
rect 664 550 694 634
rect 752 550 782 634
<< ndiff >>
rect 36 260 94 285
rect 36 226 48 260
rect 82 226 94 260
rect 36 201 94 226
rect 124 260 182 285
rect 124 226 136 260
rect 170 226 182 260
rect 124 201 182 226
rect 212 260 270 285
rect 212 226 224 260
rect 258 226 270 260
rect 212 201 270 226
rect 342 260 400 285
rect 342 226 354 260
rect 388 226 400 260
rect 342 201 400 226
rect 430 260 488 285
rect 430 226 442 260
rect 476 226 488 260
rect 430 201 488 226
rect 518 260 576 285
rect 518 226 530 260
rect 564 226 576 260
rect 518 201 576 226
rect 606 260 664 285
rect 606 226 618 260
rect 652 226 664 260
rect 606 201 664 226
rect 694 260 752 285
rect 694 226 706 260
rect 740 226 752 260
rect 694 201 752 226
rect 782 260 840 285
rect 782 226 794 260
rect 828 226 840 260
rect 782 201 840 226
<< pdiff >>
rect 36 609 94 634
rect 36 575 48 609
rect 82 575 94 609
rect 36 550 94 575
rect 124 609 182 634
rect 124 575 136 609
rect 170 575 182 609
rect 124 550 182 575
rect 212 609 270 634
rect 212 575 224 609
rect 258 575 270 609
rect 212 550 270 575
rect 342 609 400 634
rect 342 575 354 609
rect 388 575 400 609
rect 342 550 400 575
rect 430 609 488 634
rect 430 575 442 609
rect 476 575 488 609
rect 430 550 488 575
rect 518 609 576 634
rect 518 575 530 609
rect 564 575 576 609
rect 518 550 576 575
rect 606 609 664 634
rect 606 575 618 609
rect 652 575 664 609
rect 606 550 664 575
rect 694 609 752 634
rect 694 575 706 609
rect 740 575 752 609
rect 694 550 752 575
rect 782 609 840 634
rect 782 575 794 609
rect 828 575 840 609
rect 782 550 840 575
<< ndiffc >>
rect 48 226 82 260
rect 136 226 170 260
rect 224 226 258 260
rect 354 226 388 260
rect 442 226 476 260
rect 530 226 564 260
rect 618 226 652 260
rect 706 226 740 260
rect 794 226 828 260
<< pdiffc >>
rect 48 575 82 609
rect 136 575 170 609
rect 224 575 258 609
rect 354 575 388 609
rect 442 575 476 609
rect 530 575 564 609
rect 618 575 652 609
rect 706 575 740 609
rect 794 575 828 609
<< poly >>
rect 94 634 124 660
rect 182 634 212 660
rect 400 634 430 660
rect 488 634 518 660
rect 576 634 606 660
rect 664 634 694 660
rect 752 634 782 660
rect 94 518 124 550
rect 44 502 124 518
rect 44 468 60 502
rect 94 468 124 502
rect 44 452 124 468
rect 94 285 124 452
rect 182 373 212 550
rect 400 462 430 550
rect 347 444 430 462
rect 488 444 518 550
rect 576 444 606 550
rect 664 444 694 550
rect 752 444 782 550
rect 347 410 357 444
rect 391 410 782 444
rect 347 394 430 410
rect 182 357 262 373
rect 182 323 212 357
rect 246 323 262 357
rect 182 307 262 323
rect 182 285 212 307
rect 400 285 430 394
rect 488 285 518 410
rect 576 285 606 410
rect 664 285 694 410
rect 752 285 782 410
rect 94 175 124 201
rect 182 175 212 201
rect 400 175 430 201
rect 488 175 518 201
rect 576 175 606 201
rect 664 175 694 201
rect 752 175 782 201
<< polycont >>
rect 60 468 94 502
rect 357 410 391 444
rect 212 323 246 357
<< locali >>
rect 48 609 82 638
rect 48 546 82 575
rect 136 609 170 638
rect 136 546 170 575
rect 224 609 258 638
rect 224 546 258 575
rect 354 609 388 638
rect 354 546 388 575
rect 442 609 476 638
rect 44 468 60 502
rect 94 468 110 502
rect 442 496 476 575
rect 530 609 564 638
rect 530 546 564 575
rect 618 609 652 638
rect 618 496 652 575
rect 706 609 740 638
rect 706 546 740 575
rect 794 609 828 638
rect 794 496 828 575
rect 442 461 828 496
rect 794 444 828 461
rect 340 410 357 444
rect 391 410 407 444
rect 794 358 828 410
rect 48 323 60 357
rect 94 323 212 357
rect 246 323 262 357
rect 442 323 828 358
rect 48 260 82 289
rect 48 197 82 226
rect 136 260 170 289
rect 136 197 170 226
rect 224 260 258 289
rect 224 197 258 226
rect 354 260 388 289
rect 354 197 388 226
rect 442 260 476 323
rect 442 197 476 226
rect 530 260 564 289
rect 530 197 564 226
rect 618 260 652 323
rect 618 197 652 226
rect 706 260 740 289
rect 706 197 740 226
rect 794 260 828 323
rect 794 197 828 226
<< viali >>
rect 48 575 82 609
rect 136 575 170 609
rect 224 575 258 609
rect 354 575 388 609
rect 442 575 476 609
rect 60 468 94 502
rect 530 575 564 609
rect 618 575 652 609
rect 706 575 740 609
rect 794 575 828 609
rect 357 410 391 444
rect 794 410 828 444
rect 60 323 94 357
rect 48 226 82 260
rect 136 226 170 260
rect 224 226 258 260
rect 354 226 388 260
rect 442 226 476 260
rect 530 226 564 260
rect 618 226 652 260
rect 706 226 740 260
rect 794 226 828 260
<< metal1 >>
rect 0 662 876 696
rect 48 634 82 662
rect 224 634 258 662
rect 354 634 388 662
rect 530 634 564 662
rect 706 634 740 662
rect 42 609 88 634
rect 42 575 48 609
rect 82 575 88 609
rect 42 550 88 575
rect 130 609 176 634
rect 130 575 136 609
rect 170 575 176 609
rect 130 550 176 575
rect 218 609 264 634
rect 218 575 224 609
rect 258 575 264 609
rect 218 550 264 575
rect 348 609 394 634
rect 348 575 354 609
rect 388 575 394 609
rect 348 550 394 575
rect 436 609 482 634
rect 436 575 442 609
rect 476 575 482 609
rect 436 550 482 575
rect 524 609 570 634
rect 524 575 530 609
rect 564 575 570 609
rect 524 550 570 575
rect 612 609 658 634
rect 612 575 618 609
rect 652 575 658 609
rect 612 550 658 575
rect 700 609 746 634
rect 700 575 706 609
rect 740 575 746 609
rect 700 550 746 575
rect 788 609 834 634
rect 788 575 794 609
rect 828 575 834 609
rect 788 550 834 575
rect 48 502 106 508
rect 0 468 60 502
rect 94 468 106 502
rect 0 462 106 468
rect 0 410 34 462
rect 136 444 170 550
rect 345 444 403 450
rect 136 410 357 444
rect 391 410 403 444
rect 35 314 45 366
rect 97 314 107 366
rect 224 285 258 410
rect 345 404 403 410
rect 782 444 840 450
rect 782 410 794 444
rect 828 410 876 444
rect 782 404 840 410
rect 42 260 88 285
rect 42 226 48 260
rect 82 226 88 260
rect 42 201 88 226
rect 130 260 176 285
rect 130 226 136 260
rect 170 226 176 260
rect 130 201 176 226
rect 218 260 264 285
rect 218 226 224 260
rect 258 226 264 260
rect 218 201 264 226
rect 348 260 394 285
rect 348 226 354 260
rect 388 226 394 260
rect 348 201 394 226
rect 436 260 482 285
rect 436 226 442 260
rect 476 226 482 260
rect 436 201 482 226
rect 524 260 570 285
rect 524 226 530 260
rect 564 226 570 260
rect 524 201 570 226
rect 612 260 658 285
rect 612 226 618 260
rect 652 226 658 260
rect 612 201 658 226
rect 700 260 746 285
rect 700 226 706 260
rect 740 226 746 260
rect 700 201 746 226
rect 788 260 834 285
rect 788 226 794 260
rect 828 226 834 260
rect 788 201 834 226
rect 48 172 82 201
rect 354 172 388 201
rect 530 172 564 201
rect 706 172 740 201
rect 0 138 876 172
<< via1 >>
rect 45 357 97 366
rect 45 323 60 357
rect 60 323 94 357
rect 94 323 97 357
rect 45 314 97 323
<< metal2 >>
rect 45 366 97 696
rect 45 0 97 314
<< labels >>
flabel metal1 s 0 662 34 696 0 FreeSans 44 0 0 0 VDD
port 1 nsew
flabel metal1 s 0 410 34 444 0 FreeSans 44 0 0 0 A
port 2 nsew
flabel metal1 s 0 138 34 172 0 FreeSans 44 0 0 0 VSS
port 3 nsew
flabel metal2 s 45 0 97 52 0 FreeSans 44 0 0 0 WLEN
port 4 nsew
flabel metal1 s 842 410 876 444 0 FreeSans 44 0 0 0 B
port 5 nsew
<< end >>
