magic
tech sky130A
magscale 1 2
timestamp 1702731703
<< nwell >>
rect 0 2686 436 3210
rect 0 0 208 2686
<< nmos >>
rect 94 3278 124 3678
rect 312 3278 342 3678
rect 402 2432 486 2462
rect 402 2214 486 2244
rect 402 2126 486 2156
rect 404 1812 488 1842
rect 402 1504 486 1534
rect 401 1286 485 1316
rect 401 1198 485 1228
rect 411 920 495 950
rect 411 702 495 732
rect 411 614 495 644
rect 411 285 495 315
rect 411 197 495 227
<< pmos >>
rect 94 2748 124 3148
rect 312 2748 342 3148
rect 62 2432 146 2462
rect 62 2214 146 2244
rect 62 2126 146 2156
rect 62 1812 146 1842
rect 62 1504 146 1534
rect 62 1286 146 1316
rect 62 1198 146 1228
rect 62 920 146 950
rect 62 702 146 732
rect 62 614 146 644
rect 62 285 146 315
rect 62 197 146 227
<< ndiff >>
rect 36 3666 94 3678
rect 36 3290 48 3666
rect 82 3290 94 3666
rect 36 3278 94 3290
rect 124 3666 182 3678
rect 124 3290 136 3666
rect 170 3290 182 3666
rect 124 3278 182 3290
rect 254 3666 312 3678
rect 254 3290 266 3666
rect 300 3290 312 3666
rect 254 3278 312 3290
rect 342 3666 400 3678
rect 342 3290 354 3666
rect 388 3290 400 3666
rect 342 3278 400 3290
rect 402 2508 486 2520
rect 402 2474 414 2508
rect 474 2474 486 2508
rect 402 2462 486 2474
rect 402 2420 486 2432
rect 402 2386 414 2420
rect 474 2386 486 2420
rect 402 2374 486 2386
rect 402 2290 486 2302
rect 402 2256 414 2290
rect 474 2256 486 2290
rect 402 2244 486 2256
rect 402 2202 486 2214
rect 402 2168 414 2202
rect 474 2168 486 2202
rect 402 2156 486 2168
rect 402 2114 486 2126
rect 402 2080 414 2114
rect 474 2080 486 2114
rect 402 2068 486 2080
rect 404 1888 488 1900
rect 404 1854 416 1888
rect 476 1854 488 1888
rect 404 1842 488 1854
rect 404 1800 488 1812
rect 404 1766 416 1800
rect 476 1766 488 1800
rect 404 1754 488 1766
rect 402 1580 486 1592
rect 402 1546 414 1580
rect 474 1546 486 1580
rect 402 1534 486 1546
rect 402 1492 486 1504
rect 402 1458 414 1492
rect 474 1458 486 1492
rect 402 1446 486 1458
rect 401 1362 485 1374
rect 401 1328 413 1362
rect 473 1328 485 1362
rect 401 1316 485 1328
rect 401 1274 485 1286
rect 401 1240 413 1274
rect 473 1240 485 1274
rect 401 1228 485 1240
rect 401 1186 485 1198
rect 401 1152 413 1186
rect 473 1152 485 1186
rect 401 1140 485 1152
rect 411 996 495 1008
rect 411 962 423 996
rect 483 962 495 996
rect 411 950 495 962
rect 411 908 495 920
rect 411 874 423 908
rect 483 874 495 908
rect 411 862 495 874
rect 411 778 495 790
rect 411 744 423 778
rect 483 744 495 778
rect 411 732 495 744
rect 411 690 495 702
rect 411 656 423 690
rect 483 656 495 690
rect 411 644 495 656
rect 411 602 495 614
rect 411 568 423 602
rect 483 568 495 602
rect 411 556 495 568
rect 411 361 495 373
rect 411 327 423 361
rect 483 327 495 361
rect 411 315 495 327
rect 411 273 495 285
rect 411 239 423 273
rect 483 239 495 273
rect 411 227 495 239
rect 411 185 495 197
rect 411 151 423 185
rect 483 151 495 185
rect 411 139 495 151
<< pdiff >>
rect 36 3136 94 3148
rect 36 2760 48 3136
rect 82 2760 94 3136
rect 36 2748 94 2760
rect 124 3136 182 3148
rect 124 2760 136 3136
rect 170 2760 182 3136
rect 124 2748 182 2760
rect 254 3136 312 3148
rect 254 2760 266 3136
rect 300 2760 312 3136
rect 254 2748 312 2760
rect 342 3136 400 3148
rect 342 2760 354 3136
rect 388 2760 400 3136
rect 342 2748 400 2760
rect 62 2508 146 2520
rect 62 2474 74 2508
rect 134 2474 146 2508
rect 62 2462 146 2474
rect 62 2420 146 2432
rect 62 2386 74 2420
rect 134 2386 146 2420
rect 62 2374 146 2386
rect 62 2290 146 2302
rect 62 2256 74 2290
rect 134 2256 146 2290
rect 62 2244 146 2256
rect 62 2202 146 2214
rect 62 2168 74 2202
rect 134 2168 146 2202
rect 62 2156 146 2168
rect 62 2114 146 2126
rect 62 2080 74 2114
rect 134 2080 146 2114
rect 62 2068 146 2080
rect 62 1888 146 1900
rect 62 1854 74 1888
rect 134 1854 146 1888
rect 62 1842 146 1854
rect 62 1800 146 1812
rect 62 1766 74 1800
rect 134 1766 146 1800
rect 62 1754 146 1766
rect 62 1580 146 1592
rect 62 1546 74 1580
rect 134 1546 146 1580
rect 62 1534 146 1546
rect 62 1492 146 1504
rect 62 1458 74 1492
rect 134 1458 146 1492
rect 62 1446 146 1458
rect 62 1362 146 1374
rect 62 1328 74 1362
rect 134 1328 146 1362
rect 62 1316 146 1328
rect 62 1274 146 1286
rect 62 1240 74 1274
rect 134 1240 146 1274
rect 62 1228 146 1240
rect 62 1186 146 1198
rect 62 1152 74 1186
rect 134 1152 146 1186
rect 62 1140 146 1152
rect 62 996 146 1008
rect 62 962 74 996
rect 134 962 146 996
rect 62 950 146 962
rect 62 908 146 920
rect 62 874 74 908
rect 134 874 146 908
rect 62 862 146 874
rect 62 778 146 790
rect 62 744 74 778
rect 134 744 146 778
rect 62 732 146 744
rect 62 690 146 702
rect 62 656 74 690
rect 134 656 146 690
rect 62 644 146 656
rect 62 602 146 614
rect 62 568 74 602
rect 134 568 146 602
rect 62 556 146 568
rect 62 361 146 373
rect 62 327 74 361
rect 134 327 146 361
rect 62 315 146 327
rect 62 273 146 285
rect 62 239 74 273
rect 134 239 146 273
rect 62 227 146 239
rect 62 185 146 197
rect 62 151 74 185
rect 134 151 146 185
rect 62 139 146 151
<< ndiffc >>
rect 48 3290 82 3666
rect 136 3290 170 3666
rect 266 3290 300 3666
rect 354 3290 388 3666
rect 414 2474 474 2508
rect 414 2386 474 2420
rect 414 2256 474 2290
rect 414 2168 474 2202
rect 414 2080 474 2114
rect 416 1854 476 1888
rect 416 1766 476 1800
rect 414 1546 474 1580
rect 414 1458 474 1492
rect 413 1328 473 1362
rect 413 1240 473 1274
rect 413 1152 473 1186
rect 423 962 483 996
rect 423 874 483 908
rect 423 744 483 778
rect 423 656 483 690
rect 423 568 483 602
rect 423 327 483 361
rect 423 239 483 273
rect 423 151 483 185
<< pdiffc >>
rect 48 2760 82 3136
rect 136 2760 170 3136
rect 266 2760 300 3136
rect 354 2760 388 3136
rect 74 2474 134 2508
rect 74 2386 134 2420
rect 74 2256 134 2290
rect 74 2168 134 2202
rect 74 2080 134 2114
rect 74 1854 134 1888
rect 74 1766 134 1800
rect 74 1546 134 1580
rect 74 1458 134 1492
rect 74 1328 134 1362
rect 74 1240 134 1274
rect 74 1152 134 1186
rect 74 962 134 996
rect 74 874 134 908
rect 74 744 134 778
rect 74 656 134 690
rect 74 568 134 602
rect 74 327 134 361
rect 74 239 134 273
rect 74 151 134 185
<< psubdiff >>
rect 420 473 528 485
rect 420 439 444 473
rect 504 439 528 473
rect 420 427 528 439
<< nsubdiff >>
rect 50 488 158 500
rect 50 454 74 488
rect 134 454 158 488
rect 50 442 158 454
<< psubdiffcont >>
rect 444 439 504 473
<< nsubdiffcont >>
rect 74 454 134 488
<< poly >>
rect 94 3678 124 3704
rect 312 3678 342 3704
rect 94 3148 124 3278
rect 193 3230 260 3247
rect 312 3230 342 3278
rect 193 3195 209 3230
rect 243 3195 342 3230
rect 193 3179 260 3195
rect 312 3148 342 3195
rect 94 2702 124 2748
rect 312 2722 342 2748
rect 94 2686 174 2702
rect 94 2652 124 2686
rect 158 2652 174 2686
rect 94 2636 174 2652
rect 184 2496 250 2512
rect 184 2462 200 2496
rect 234 2462 250 2496
rect 36 2432 62 2462
rect 146 2432 250 2462
rect 296 2496 362 2512
rect 296 2462 312 2496
rect 346 2462 362 2496
rect 296 2432 402 2462
rect 486 2432 512 2462
rect 207 2278 274 2294
rect 207 2244 223 2278
rect 258 2244 274 2278
rect 36 2214 62 2244
rect 146 2214 402 2244
rect 486 2214 512 2244
rect 36 2126 62 2156
rect 146 2126 402 2156
rect 486 2126 512 2156
rect 223 2042 258 2126
rect 207 2026 274 2042
rect 207 1992 223 2026
rect 258 1992 274 2026
rect 207 1976 274 1992
rect 320 1958 386 1974
rect 320 1924 336 1958
rect 370 1924 386 1958
rect 320 1908 386 1924
rect 194 1876 260 1892
rect 194 1842 210 1876
rect 244 1842 260 1876
rect 36 1812 62 1842
rect 146 1812 260 1842
rect 348 1842 378 1908
rect 348 1812 404 1842
rect 488 1812 514 1842
rect 320 1650 386 1666
rect 320 1616 336 1650
rect 370 1616 386 1650
rect 320 1600 386 1616
rect 194 1568 260 1584
rect 194 1534 210 1568
rect 244 1534 260 1568
rect 36 1504 62 1534
rect 146 1504 260 1534
rect 356 1534 386 1600
rect 356 1504 402 1534
rect 486 1504 512 1534
rect 194 1350 260 1366
rect 194 1316 210 1350
rect 244 1316 260 1350
rect 36 1286 62 1316
rect 146 1286 401 1316
rect 485 1286 511 1316
rect 36 1198 62 1228
rect 146 1198 401 1228
rect 485 1198 511 1228
rect 261 1112 295 1198
rect 245 1096 311 1112
rect 245 1062 261 1096
rect 295 1062 311 1096
rect 245 1046 311 1062
rect 184 984 250 1000
rect 184 950 200 984
rect 234 950 250 984
rect 36 920 62 950
rect 146 920 250 950
rect 306 984 373 1001
rect 306 950 322 984
rect 356 950 373 984
rect 306 920 411 950
rect 495 920 521 950
rect 323 766 389 782
rect 323 732 339 766
rect 373 732 389 766
rect 36 702 62 732
rect 146 702 411 732
rect 495 702 521 732
rect 36 614 62 644
rect 146 614 411 644
rect 495 614 521 644
rect 339 533 373 614
rect 323 517 389 533
rect 323 483 339 517
rect 373 483 389 517
rect 323 467 389 483
rect 192 349 258 365
rect 192 315 208 349
rect 242 315 258 349
rect 36 285 62 315
rect 146 285 411 315
rect 495 285 521 315
rect 36 197 62 227
rect 146 197 411 227
rect 495 197 521 227
rect 208 111 242 197
rect 192 101 258 111
rect 192 67 208 101
rect 242 67 258 101
rect 192 51 258 67
<< polycont >>
rect 209 3195 243 3230
rect 124 2652 158 2686
rect 200 2462 234 2496
rect 312 2462 346 2496
rect 223 2244 258 2278
rect 223 1992 258 2026
rect 336 1924 370 1958
rect 210 1842 244 1876
rect 336 1616 370 1650
rect 210 1534 244 1568
rect 210 1316 244 1350
rect 261 1062 295 1096
rect 200 950 234 984
rect 322 950 356 984
rect 339 732 373 766
rect 339 483 373 517
rect 208 315 242 349
rect 208 67 242 101
<< locali >>
rect 48 3666 82 3682
rect 48 3274 82 3290
rect 136 3666 170 3682
rect 136 3230 170 3290
rect 266 3666 300 3682
rect 266 3274 300 3290
rect 354 3666 388 3682
rect 354 3274 388 3290
rect 136 3195 209 3230
rect 243 3195 260 3230
rect 48 3136 82 3152
rect 48 2744 82 2760
rect 136 3136 170 3195
rect 136 2744 170 2760
rect 266 3136 300 3152
rect 266 2744 300 2760
rect 354 3136 388 3152
rect 354 2744 388 2760
rect 108 2652 124 2686
rect 158 2652 174 2686
rect 116 2535 433 2569
rect 116 2508 150 2535
rect 58 2474 74 2508
rect 134 2474 150 2508
rect 398 2508 433 2535
rect 184 2462 200 2496
rect 234 2462 250 2496
rect 296 2462 312 2496
rect 346 2462 362 2496
rect 398 2474 414 2508
rect 474 2474 558 2508
rect 58 2386 74 2420
rect 134 2386 414 2420
rect 474 2386 490 2420
rect 87 2290 121 2386
rect 58 2256 74 2290
rect 134 2256 150 2290
rect 223 2278 258 2294
rect 428 2290 462 2386
rect 398 2256 414 2290
rect 474 2256 490 2290
rect 58 2168 74 2202
rect 134 2168 150 2202
rect 223 2114 258 2244
rect 398 2168 414 2202
rect 474 2168 490 2202
rect 58 2080 74 2114
rect 134 2080 257 2114
rect 291 2080 414 2114
rect 474 2080 490 2114
rect 524 2026 558 2474
rect 86 1992 223 2026
rect 258 1992 558 2026
rect 86 1888 120 1992
rect 208 1924 336 1958
rect 370 1924 386 1958
rect 438 1888 472 1992
rect 58 1854 74 1888
rect 134 1854 150 1888
rect 194 1842 210 1876
rect 244 1842 331 1876
rect 400 1854 416 1888
rect 476 1854 492 1888
rect 58 1766 74 1800
rect 134 1766 416 1800
rect 476 1766 558 1800
rect 86 1684 261 1718
rect 295 1684 472 1718
rect 86 1580 120 1684
rect 208 1616 336 1650
rect 370 1616 386 1650
rect 438 1580 472 1684
rect 58 1546 74 1580
rect 134 1546 150 1580
rect 194 1534 210 1568
rect 244 1534 330 1568
rect 398 1546 414 1580
rect 474 1546 490 1580
rect 58 1458 74 1492
rect 134 1458 414 1492
rect 474 1458 490 1492
rect 86 1362 120 1458
rect 58 1328 74 1362
rect 134 1328 150 1362
rect 210 1350 244 1366
rect 435 1362 469 1458
rect 397 1328 413 1362
rect 473 1328 489 1362
rect 58 1240 74 1274
rect 134 1240 150 1274
rect 210 1186 244 1316
rect 397 1240 413 1274
rect 473 1240 489 1274
rect 524 1186 558 1766
rect 58 1152 74 1186
rect 134 1152 413 1186
rect 473 1152 558 1186
rect 116 1062 261 1096
rect 295 1062 441 1096
rect 116 996 150 1062
rect 58 962 74 996
rect 134 962 150 996
rect 407 996 441 1062
rect 184 950 200 984
rect 234 950 250 984
rect 306 950 322 984
rect 356 950 373 984
rect 407 962 423 996
rect 483 962 499 996
rect 58 874 74 908
rect 134 874 423 908
rect 483 874 499 908
rect 86 778 120 874
rect 58 744 74 778
rect 134 744 150 778
rect 339 766 373 782
rect 435 778 469 874
rect 407 744 423 778
rect 483 744 499 778
rect 58 656 74 690
rect 134 656 150 690
rect 339 602 373 732
rect 407 656 423 690
rect 483 656 499 690
rect 58 568 74 602
rect 134 568 423 602
rect 483 568 499 602
rect 339 517 373 533
rect 58 454 74 488
rect 134 454 150 488
rect 208 413 261 447
rect 58 327 74 361
rect 134 327 150 361
rect 208 349 242 413
rect 58 239 74 273
rect 134 239 150 273
rect 208 185 242 315
rect 339 273 373 483
rect 428 439 444 473
rect 504 439 520 473
rect 407 327 423 361
rect 483 327 499 361
rect 407 239 423 273
rect 483 239 499 273
rect 58 151 74 185
rect 134 151 423 185
rect 483 151 499 185
rect 208 101 242 117
rect 208 51 242 67
<< viali >>
rect 48 3290 82 3666
rect 136 3290 170 3666
rect 266 3290 300 3666
rect 354 3290 388 3666
rect 48 2760 82 3136
rect 136 2760 170 3136
rect 266 2760 300 3136
rect 354 2760 388 3136
rect 124 2652 158 2686
rect 74 2474 134 2508
rect 200 2462 234 2496
rect 312 2462 346 2496
rect 414 2474 474 2508
rect 74 2386 134 2420
rect 414 2386 474 2420
rect 74 2256 134 2290
rect 414 2256 474 2290
rect 74 2168 134 2202
rect 414 2168 474 2202
rect 74 2080 134 2114
rect 257 2080 291 2114
rect 414 2080 474 2114
rect 174 1924 208 1958
rect 74 1854 134 1888
rect 331 1842 365 1876
rect 416 1854 476 1888
rect 74 1766 134 1800
rect 416 1766 476 1800
rect 261 1684 295 1718
rect 174 1616 208 1650
rect 74 1546 134 1580
rect 330 1534 364 1568
rect 414 1546 474 1580
rect 74 1458 134 1492
rect 414 1458 474 1492
rect 74 1328 134 1362
rect 413 1328 473 1362
rect 74 1240 134 1274
rect 413 1240 473 1274
rect 74 1152 134 1186
rect 413 1152 473 1186
rect 261 1062 295 1096
rect 74 962 134 996
rect 200 950 234 984
rect 322 950 356 984
rect 423 962 483 996
rect 74 874 134 908
rect 423 874 483 908
rect 74 744 134 778
rect 423 744 483 778
rect 74 656 134 690
rect 423 656 483 690
rect 74 568 134 602
rect 423 568 483 602
rect 87 454 121 488
rect 261 413 295 447
rect 74 327 134 361
rect 74 239 134 273
rect 457 439 491 473
rect 423 327 483 361
rect 339 239 373 273
rect 423 239 483 273
rect 74 151 134 185
rect 423 151 483 185
rect 208 67 242 101
<< metal1 >>
rect 463 3861 497 3901
rect 463 3827 612 3861
rect 48 3758 469 3792
rect 48 3678 82 3758
rect 117 3678 127 3730
rect 179 3678 189 3730
rect 266 3678 300 3758
rect 335 3678 345 3730
rect 397 3678 407 3730
rect 42 3666 88 3678
rect 42 3290 48 3666
rect 82 3290 88 3666
rect 42 3278 88 3290
rect 130 3666 176 3678
rect 130 3290 136 3666
rect 170 3290 176 3666
rect 130 3278 176 3290
rect 260 3666 306 3678
rect 260 3290 266 3666
rect 300 3290 306 3666
rect 260 3278 306 3290
rect 348 3666 394 3678
rect 348 3290 354 3666
rect 388 3290 394 3666
rect 348 3278 394 3290
rect 47 3176 301 3210
rect 47 3148 82 3176
rect 266 3148 301 3176
rect 354 3148 388 3278
rect 435 3225 469 3758
rect 578 3566 612 3827
rect 568 3514 578 3566
rect 630 3514 640 3566
rect 435 3191 559 3225
rect 42 3136 88 3148
rect 42 2760 48 3136
rect 82 2760 88 3136
rect 42 2748 88 2760
rect 130 3136 176 3148
rect 130 2760 136 3136
rect 170 2760 176 3136
rect 130 2748 176 2760
rect 260 3136 306 3148
rect 260 2760 266 3136
rect 300 2760 306 3136
rect 260 2748 306 2760
rect 348 3136 394 3148
rect 348 2760 354 3136
rect 388 2760 394 3136
rect 348 2748 394 2760
rect 47 2720 82 2748
rect 0 2686 82 2720
rect 112 2686 170 2692
rect 525 2686 559 3191
rect 0 2202 34 2686
rect 112 2652 124 2686
rect 158 2652 286 2686
rect 112 2646 170 2652
rect 244 2631 286 2652
rect 244 2621 296 2631
rect 244 2559 296 2569
rect 62 2508 146 2514
rect 402 2508 486 2514
rect 62 2474 74 2508
rect 134 2474 146 2508
rect 62 2468 146 2474
rect 174 2496 240 2508
rect 174 2462 200 2496
rect 234 2462 240 2496
rect 174 2450 240 2462
rect 304 2496 373 2508
rect 304 2462 312 2496
rect 346 2462 373 2496
rect 402 2474 414 2508
rect 474 2474 486 2508
rect 402 2468 486 2474
rect 62 2420 146 2426
rect 62 2386 74 2420
rect 134 2386 146 2420
rect 62 2380 146 2386
rect 62 2290 146 2296
rect 62 2256 74 2290
rect 134 2256 146 2290
rect 62 2250 146 2256
rect 62 2202 146 2208
rect 0 2168 74 2202
rect 134 2168 146 2202
rect 0 1274 34 2168
rect 62 2162 146 2168
rect 62 2114 146 2120
rect 62 2080 74 2114
rect 134 2080 146 2114
rect 62 2074 146 2080
rect 174 1970 208 2450
rect 304 2449 373 2462
rect 248 2123 300 2133
rect 248 2061 300 2071
rect 168 1958 214 1970
rect 168 1924 174 1958
rect 208 1924 214 1958
rect 168 1912 214 1924
rect 62 1888 146 1894
rect 62 1854 74 1888
rect 134 1854 146 1888
rect 62 1848 146 1854
rect 62 1800 146 1806
rect 62 1766 74 1800
rect 134 1766 146 1800
rect 62 1760 146 1766
rect 174 1662 208 1912
rect 339 1888 373 2449
rect 402 2420 486 2426
rect 402 2386 414 2420
rect 474 2386 486 2420
rect 402 2380 486 2386
rect 525 2364 558 2686
rect 402 2290 486 2296
rect 402 2256 414 2290
rect 474 2256 486 2290
rect 402 2250 486 2256
rect 402 2202 486 2208
rect 524 2202 558 2364
rect 402 2168 414 2202
rect 474 2168 558 2202
rect 402 2162 486 2168
rect 402 2114 486 2120
rect 402 2080 414 2114
rect 474 2080 486 2114
rect 402 2074 486 2080
rect 524 1921 558 2168
rect 325 1876 373 1888
rect 325 1842 331 1876
rect 365 1842 373 1876
rect 404 1888 488 1894
rect 404 1854 416 1888
rect 476 1854 488 1888
rect 404 1848 488 1854
rect 325 1830 373 1842
rect 255 1718 301 1730
rect 255 1684 261 1718
rect 295 1684 301 1718
rect 255 1672 301 1684
rect 168 1650 214 1662
rect 168 1616 174 1650
rect 208 1616 214 1650
rect 168 1604 214 1616
rect 62 1580 146 1586
rect 62 1546 74 1580
rect 134 1546 146 1580
rect 62 1540 146 1546
rect 62 1492 146 1498
rect 62 1458 74 1492
rect 134 1458 146 1492
rect 62 1452 146 1458
rect 62 1362 146 1368
rect 62 1328 74 1362
rect 134 1328 146 1362
rect 62 1322 146 1328
rect 62 1274 146 1280
rect 0 1240 74 1274
rect 134 1240 146 1274
rect 0 690 34 1240
rect 62 1234 146 1240
rect 62 1186 146 1192
rect 62 1152 74 1186
rect 134 1152 146 1186
rect 62 1146 146 1152
rect 62 996 146 1002
rect 62 962 74 996
rect 134 962 146 996
rect 62 956 146 962
rect 174 996 208 1604
rect 261 1108 295 1672
rect 339 1580 373 1830
rect 404 1800 488 1806
rect 404 1766 416 1800
rect 476 1766 488 1800
rect 404 1760 488 1766
rect 324 1568 373 1580
rect 324 1534 330 1568
rect 364 1534 373 1568
rect 402 1580 486 1586
rect 402 1546 414 1580
rect 474 1546 486 1580
rect 402 1540 486 1546
rect 324 1522 373 1534
rect 255 1096 301 1108
rect 255 1062 261 1096
rect 295 1062 301 1096
rect 255 1050 301 1062
rect 339 996 373 1522
rect 402 1492 486 1498
rect 402 1458 414 1492
rect 474 1458 486 1492
rect 402 1452 486 1458
rect 401 1362 485 1368
rect 401 1328 413 1362
rect 473 1328 485 1362
rect 401 1322 485 1328
rect 401 1274 485 1280
rect 525 1274 558 1921
rect 401 1240 413 1274
rect 473 1240 558 1274
rect 401 1234 485 1240
rect 401 1186 485 1192
rect 401 1152 413 1186
rect 473 1152 485 1186
rect 401 1146 485 1152
rect 174 984 240 996
rect 174 950 200 984
rect 234 950 240 984
rect 174 938 240 950
rect 316 984 373 996
rect 316 950 322 984
rect 356 950 373 984
rect 411 996 495 1002
rect 411 962 423 996
rect 483 962 495 996
rect 411 956 495 962
rect 316 938 373 950
rect 62 908 146 914
rect 62 874 74 908
rect 134 874 146 908
rect 62 868 146 874
rect 62 778 146 784
rect 62 744 74 778
rect 134 744 146 778
rect 62 738 146 744
rect 62 690 146 696
rect 0 656 74 690
rect 134 656 146 690
rect 0 488 34 656
rect 62 650 146 656
rect 62 602 146 608
rect 62 568 74 602
rect 134 568 146 602
rect 62 562 146 568
rect 81 488 127 500
rect 0 454 87 488
rect 121 454 127 488
rect 0 273 34 454
rect 81 442 127 454
rect 62 361 146 367
rect 174 361 208 938
rect 255 447 301 459
rect 339 447 373 938
rect 411 908 495 914
rect 411 874 423 908
rect 483 874 495 908
rect 411 868 495 874
rect 411 778 495 784
rect 411 744 423 778
rect 483 744 495 778
rect 411 738 495 744
rect 411 690 495 696
rect 524 690 558 1240
rect 411 656 423 690
rect 483 656 558 690
rect 411 650 495 656
rect 411 602 495 608
rect 411 568 423 602
rect 483 568 495 602
rect 411 562 495 568
rect 524 485 558 656
rect 255 413 261 447
rect 295 413 373 447
rect 451 473 558 485
rect 451 439 457 473
rect 491 439 558 473
rect 451 427 558 439
rect 255 401 301 413
rect 411 361 495 367
rect 62 327 74 361
rect 134 327 423 361
rect 483 327 495 361
rect 62 321 146 327
rect 411 321 495 327
rect 62 273 146 279
rect 0 239 74 273
rect 134 239 146 273
rect 0 0 34 239
rect 62 233 146 239
rect 333 273 379 285
rect 333 239 339 273
rect 373 239 379 273
rect 333 227 379 239
rect 411 273 495 279
rect 524 273 558 427
rect 411 239 423 273
rect 483 239 558 273
rect 411 233 495 239
rect 62 185 146 191
rect 62 151 74 185
rect 134 151 146 185
rect 62 145 146 151
rect 202 101 248 113
rect 202 67 208 101
rect 242 67 248 101
rect 202 55 248 67
rect 208 0 242 55
rect 339 0 373 227
rect 411 185 495 191
rect 411 151 423 185
rect 483 151 495 185
rect 411 145 495 151
rect 524 0 558 239
rect 620 85 630 137
rect 682 85 692 137
rect 620 0 654 85
<< via1 >>
rect 127 3678 179 3730
rect 345 3678 397 3730
rect 578 3514 630 3566
rect 244 2569 296 2621
rect 248 2114 300 2123
rect 248 2080 257 2114
rect 257 2080 291 2114
rect 291 2080 300 2114
rect 248 2071 300 2080
rect 630 85 682 137
<< metal2 >>
rect 164 3740 216 3901
rect 127 3730 219 3740
rect 179 3678 219 3730
rect 127 3668 219 3678
rect 345 3730 397 3740
rect 488 3730 540 3901
rect 397 3678 540 3730
rect 345 3668 397 3678
rect 578 3566 630 3576
rect 630 3514 772 3566
rect 578 3507 630 3514
rect 234 2569 244 2621
rect 296 2569 306 2621
rect 253 2123 287 2569
rect 238 2071 248 2123
rect 300 2071 310 2123
rect 630 137 682 147
rect 720 137 772 3514
rect 682 85 772 137
rect 630 75 682 85
<< labels >>
rlabel metal2 164 3849 216 3901 0 DW_
rlabel metal2 488 3849 540 3901 0 DW
rlabel metal1 0 0 34 35 0 VDD
rlabel metal1 208 0 242 35 0 clk
rlabel metal1 339 0 373 35 0 d
rlabel metal1 524 0 558 35 0 VSS
rlabel metal1 620 0 654 35 0 SB
<< end >>
