magic
tech sky130A
magscale 1 2
timestamp 1703326108
<< nwell >>
rect 0 488 482 696
<< nmos >>
rect 94 200 124 284
rect 182 200 212 284
rect 270 200 300 284
rect 358 200 388 284
<< pmos >>
rect 94 550 124 634
rect 182 550 212 634
rect 270 550 300 634
rect 358 550 388 634
<< ndiff >>
rect 36 272 94 284
rect 36 212 48 272
rect 82 212 94 272
rect 36 200 94 212
rect 124 272 182 284
rect 124 212 136 272
rect 170 212 182 272
rect 124 200 182 212
rect 212 272 270 284
rect 212 212 224 272
rect 258 212 270 272
rect 212 200 270 212
rect 300 272 358 284
rect 300 212 312 272
rect 346 212 358 272
rect 300 200 358 212
rect 388 272 446 284
rect 388 212 400 272
rect 434 212 446 272
rect 388 200 446 212
<< pdiff >>
rect 36 622 94 634
rect 36 562 48 622
rect 82 562 94 622
rect 36 550 94 562
rect 124 622 182 634
rect 124 562 136 622
rect 170 562 182 622
rect 124 550 182 562
rect 212 622 270 634
rect 212 562 224 622
rect 258 562 270 622
rect 212 550 270 562
rect 300 622 358 634
rect 300 562 312 622
rect 346 562 358 622
rect 300 550 358 562
rect 388 622 446 634
rect 388 562 400 622
rect 434 562 446 622
rect 388 550 446 562
<< ndiffc >>
rect 48 212 82 272
rect 136 212 170 272
rect 224 212 258 272
rect 312 212 346 272
rect 400 212 434 272
<< pdiffc >>
rect 48 562 82 622
rect 136 562 170 622
rect 224 562 258 622
rect 312 562 346 622
rect 400 562 434 622
<< poly >>
rect 94 634 124 660
rect 182 634 212 660
rect 270 634 300 660
rect 358 634 388 660
rect 94 513 124 550
rect 44 503 124 513
rect 182 509 212 550
rect 44 469 60 503
rect 94 469 124 503
rect 44 459 124 469
rect 94 284 124 459
rect 170 493 225 509
rect 170 459 180 493
rect 214 459 225 493
rect 170 443 225 459
rect 182 284 212 443
rect 270 373 300 550
rect 258 357 312 373
rect 258 323 268 357
rect 302 323 312 357
rect 258 307 312 323
rect 270 284 300 307
rect 358 284 388 550
rect 94 174 124 200
rect 182 174 212 200
rect 270 174 300 200
rect 358 141 388 200
rect 346 125 400 141
rect 346 91 356 125
rect 390 91 400 125
rect 346 75 400 91
<< polycont >>
rect 60 469 94 503
rect 180 459 214 493
rect 268 323 302 357
rect 356 91 390 125
<< locali >>
rect 48 622 82 638
rect 48 546 82 562
rect 136 622 170 638
rect 136 546 170 562
rect 224 622 258 638
rect 224 546 258 562
rect 312 622 346 638
rect 312 546 346 562
rect 400 622 434 638
rect 400 546 434 562
rect 44 469 60 503
rect 94 469 110 503
rect 180 493 214 509
rect 180 429 214 459
rect 252 323 268 357
rect 302 323 318 357
rect 48 272 82 288
rect 48 196 82 212
rect 136 272 170 288
rect 136 196 170 212
rect 224 272 258 288
rect 224 196 258 212
rect 312 272 346 288
rect 312 196 346 212
rect 400 272 434 288
rect 400 196 434 212
rect 356 125 390 141
rect 356 82 390 91
<< viali >>
rect 48 562 82 622
rect 136 562 170 622
rect 224 562 258 622
rect 312 562 346 622
rect 400 562 434 622
rect 60 469 94 503
rect 180 395 214 429
rect 268 323 302 355
rect 268 321 302 323
rect 48 212 82 272
rect 136 212 170 272
rect 224 212 258 272
rect 312 212 346 272
rect 400 212 434 272
rect 356 48 390 82
<< metal1 >>
rect 0 662 482 696
rect 48 634 82 662
rect 224 634 258 662
rect 400 634 434 662
rect 42 622 88 634
rect 42 562 48 622
rect 82 562 88 622
rect 42 550 88 562
rect 130 622 176 634
rect 130 562 136 622
rect 170 562 176 622
rect 130 550 176 562
rect 218 622 264 634
rect 218 562 224 622
rect 258 562 264 622
rect 218 550 264 562
rect 306 622 352 634
rect 306 562 312 622
rect 346 562 352 622
rect 306 550 352 562
rect 394 622 440 634
rect 394 562 400 622
rect 434 562 440 622
rect 394 550 440 562
rect 136 514 170 550
rect 312 514 346 550
rect 48 503 106 509
rect 0 469 60 503
rect 94 469 106 503
rect 136 480 434 514
rect 48 463 106 469
rect 400 444 434 480
rect 168 429 226 435
rect 0 395 180 429
rect 214 395 226 429
rect 168 389 226 395
rect 400 410 482 444
rect 256 355 314 361
rect 0 321 268 355
rect 302 321 314 355
rect 256 315 314 321
rect 400 284 434 410
rect 42 272 88 284
rect 42 212 48 272
rect 82 212 88 272
rect 42 200 88 212
rect 130 272 176 284
rect 130 212 136 272
rect 170 212 176 272
rect 130 200 176 212
rect 218 272 264 284
rect 218 212 224 272
rect 258 212 264 272
rect 218 200 264 212
rect 306 272 352 284
rect 306 212 312 272
rect 346 212 352 272
rect 306 200 352 212
rect 394 272 440 284
rect 394 212 400 272
rect 434 212 440 272
rect 394 200 440 212
rect 48 172 82 200
rect 0 138 482 172
rect 344 82 402 88
rect 0 48 356 82
rect 390 48 402 82
rect 344 42 402 48
<< labels >>
rlabel metal1 0 662 34 696 0 VDD
rlabel metal1 0 469 34 503 0 A
rlabel metal1 0 395 34 429 0 B
rlabel metal1 0 321 34 355 0 C
rlabel metal1 0 138 34 172 0 VSS
rlabel metal1 0 48 34 82 0 D
rlabel metal1 448 410 482 444 0 Y
<< end >>
