magic
tech sky130A
magscale 1 2
timestamp 1703586605
<< error_s >>
rect 1344 165 1420 199
<< metal1 >>
rect 1279 509 1289 565
rect 1345 509 1355 565
rect 1279 444 1313 509
rect 1206 410 1313 444
rect 1344 165 1420 199
<< via1 >>
rect 1289 509 1345 565
<< metal2 >>
rect -149 1433 -97 1726
rect 1289 565 1345 575
rect 1289 499 1345 509
<< via2 >>
rect 1289 509 1345 565
<< metal3 >>
rect 1249 565 1420 570
rect 1249 509 1289 565
rect 1345 509 1420 565
rect 1249 504 1420 509
use not_f  not_f_0 ~/Desktop/FabRAM/FE/sram130/not
timestamp 1703586424
transform 1 0 0 0 1 0
box 0 138 330 696
use row_driver_f  row_driver_f_0 ~/Desktop/FabRAM/FE/sram130/row_driver
timestamp 1703586424
transform 1 0 330 0 1 0
box 0 0 876 696
<< end >>
