magic
tech sky130A
magscale 1 2
timestamp 1703664456
<< metal1 >>
rect 2179 606 2213 1076
rect 2179 572 2289 606
rect 1341 -651 1351 -629
rect 831 -685 1351 -651
rect 1407 -685 1417 -629
rect 1437 -1347 1447 -1325
rect 831 -1381 1447 -1347
rect 1503 -1381 1513 -1325
rect 1544 -2043 1554 -2021
rect 831 -2077 1554 -2043
rect 1610 -2077 1620 -2021
rect 1642 -2739 1652 -2717
rect 831 -2773 1652 -2739
rect 1708 -2773 1718 -2717
<< via1 >>
rect 1351 -685 1407 -629
rect 1447 -1381 1503 -1325
rect 1554 -2077 1610 -2021
rect 1652 -2773 1708 -2717
<< metal2 >>
rect 1351 1858 1407 1868
rect 1351 1792 1407 1802
rect 1351 -619 1406 1792
rect 1447 1732 1503 1742
rect 1351 -629 1407 -619
rect 1351 -695 1407 -685
rect 1447 -1325 1503 1676
rect 1447 -1394 1503 -1381
rect 1554 1606 1610 1616
rect 1554 -2021 1610 1550
rect 1554 -2087 1610 -2077
rect 1652 1480 1708 1490
rect 1652 -2717 1708 1424
rect 1652 -2783 1708 -2773
<< via2 >>
rect 1351 1802 1407 1858
rect 1447 1676 1503 1732
rect 1554 1550 1610 1606
rect 1652 1424 1708 1480
<< metal3 >>
rect 1341 1858 2289 1863
rect 1341 1802 1351 1858
rect 1407 1802 2289 1858
rect 1341 1797 2289 1802
rect 1437 1732 2289 1737
rect 1437 1676 1447 1732
rect 1503 1676 2289 1732
rect 1437 1671 2289 1676
rect 1544 1606 2289 1611
rect 1544 1550 1554 1606
rect 1610 1550 2289 1606
rect 1544 1545 2289 1550
rect 1642 1480 2289 1485
rect 1642 1424 1652 1480
rect 1708 1424 2289 1480
rect 1642 1419 2289 1424
use col_dec4_f  col_dec4_f_1
timestamp 1703662019
transform 1 0 0 0 1 0
box 0 0 2300 2492
<< end >>
