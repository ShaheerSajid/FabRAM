magic
tech sky130A
magscale 1 2
timestamp 1702483994
<< error_s >>
rect 123 14 181 20
rect 123 -20 135 14
rect 123 -26 181 -20
<< nwell >>
rect -199 0 0 324
rect 19 0 262 1
rect 306 0 521 324
rect -199 -224 -174 0
rect 44 -39 262 0
rect 44 -208 46 -39
rect 480 -224 521 0
rect -200 -962 -174 -754
rect 132 -962 174 -754
rect 480 -962 521 -754
<< psubdiff >>
rect -174 -596 -92 -577
rect -174 -656 -150 -596
rect -116 -656 -92 -596
rect -174 -685 -92 -656
<< nsubdiff >>
rect -102 139 -20 163
rect -102 79 -77 139
rect -43 79 -20 139
rect -102 55 -20 79
<< psubdiffcont >>
rect -150 -656 -116 -596
<< nsubdiffcont >>
rect -77 79 -43 139
<< poly >>
rect 94 14 212 36
rect 94 6 135 14
rect 119 -20 135 6
rect 169 6 212 14
rect 169 -20 185 6
rect 119 -36 185 -20
rect 138 -75 168 -36
rect -80 -370 -50 -188
rect 356 -350 386 -162
rect 356 -366 436 -350
rect 356 -370 386 -366
rect -80 -400 386 -370
rect 420 -400 436 -366
rect 370 -416 436 -400
rect 20 -741 386 -711
rect 286 -742 386 -741
rect 356 -790 386 -742
rect -80 -947 -50 -926
rect -156 -977 -50 -947
rect -80 -1004 -50 -977
rect 8 -938 38 -926
rect 8 -954 88 -938
rect 268 -946 298 -926
rect 8 -988 38 -954
rect 72 -988 88 -954
rect 215 -976 298 -946
rect 8 -1004 88 -988
rect 268 -1005 298 -976
rect 356 -938 386 -926
rect 356 -954 436 -938
rect 356 -988 386 -954
rect 420 -988 436 -954
rect 356 -1004 436 -988
<< polycont >>
rect 135 -20 169 14
rect 386 -400 420 -366
rect 38 -988 72 -954
rect 386 -988 420 -954
<< locali >>
rect -77 300 170 334
rect -77 155 -43 300
rect 136 266 170 300
rect -91 139 -29 155
rect -91 79 -77 139
rect -43 79 -29 139
rect -91 63 -29 79
rect 48 -92 82 58
rect 119 -20 135 14
rect 169 -20 185 14
rect 224 -92 258 58
rect 48 -126 126 -92
rect 180 -126 258 -92
rect -38 -271 -4 -166
rect 310 -271 344 -166
rect -38 -305 92 -271
rect 180 -305 344 -271
rect -26 -481 8 -305
rect 298 -481 332 -305
rect 370 -400 386 -366
rect 420 -400 436 -366
rect -166 -596 -100 -580
rect -166 -656 -150 -596
rect -116 -656 -100 -596
rect -166 -672 -100 -656
rect -150 -724 -116 -672
rect -150 -758 171 -724
rect 20 -759 171 -758
rect -126 -954 -92 -904
rect -126 -988 38 -954
rect 72 -988 88 -954
rect -126 -1026 -92 -988
rect 137 -1155 171 -759
rect 398 -812 432 -400
rect 222 -954 256 -904
rect 222 -988 386 -954
rect 420 -988 436 -954
rect 222 -1026 256 -988
rect 137 -1192 171 -1189
<< viali >>
rect 135 -20 169 14
rect 137 -1189 171 -1155
<< metal1 >>
rect -199 308 521 342
rect -171 228 -161 280
rect -109 262 -99 280
rect 136 262 170 308
rect 419 262 429 280
rect -109 228 82 262
rect 224 228 429 262
rect 481 228 491 280
rect 123 14 181 20
rect 123 -20 135 14
rect 169 -20 185 14
rect 123 -26 181 -20
rect -200 -778 521 -738
rect -38 -816 -4 -778
rect 310 -816 344 -778
rect 50 -1030 84 -900
rect 398 -1030 432 -900
rect -38 -1152 -4 -1102
rect 125 -1152 183 -1149
rect 310 -1152 344 -1102
rect -200 -1155 521 -1152
rect -200 -1189 137 -1155
rect 171 -1189 521 -1155
rect -200 -1192 521 -1189
rect 125 -1195 183 -1192
<< via1 >>
rect -161 228 -109 280
rect 429 228 481 280
<< metal2 >>
rect -161 280 -109 376
rect -161 218 -109 228
rect 429 280 481 376
rect 429 218 481 228
use sky130_fd_pr__pfet_01v8_5SMHNA  m1
timestamp 1702473764
transform -1 0 109 0 1 162
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_523TXA  m4
timestamp 1702478055
transform 1 0 -65 0 1 -112
box -109 -112 109 112
use sky130_fd_pr__pfet_01v8_523TXA  m5
timestamp 1702478055
transform -1 0 371 0 1 -112
box -109 -112 109 112
use sky130_fd_pr__nfet_01v8_L8ATA9  m6
timestamp 1702478055
transform -1 0 35 0 1 -585
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_L8ATA9  m7
timestamp 1702478055
transform 1 0 271 0 1 -585
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_A6LSUL  m8 ~/Desktop/FabRAM/FE/sram130/common
timestamp 1702483205
transform -1 0 -65 0 1 -1072
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m9 ~/Desktop/FabRAM/FE/sram130/common
timestamp 1702483205
transform -1 0 -65 0 1 -858
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m10
timestamp 1702483205
transform 1 0 23 0 1 -858
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_A6LSUL  m11
timestamp 1702483205
transform 1 0 23 0 1 -1072
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_A6LSUL  m12
timestamp 1702483205
transform -1 0 283 0 1 -1072
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m13
timestamp 1702483205
transform -1 0 283 0 1 -858
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m14
timestamp 1702483205
transform 1 0 371 0 1 -858
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_A6LSUL  m15
timestamp 1702483205
transform 1 0 371 0 1 -1072
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_5SMHNA  sky130_fd_pr__pfet_01v8_5SMHNA_0
timestamp 1702473764
transform 1 0 197 0 1 162
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_5SMHNA  sky130_fd_pr__pfet_01v8_5SMHNA_1
timestamp 1702473764
transform 1 0 153 0 1 -201
box -109 -162 109 162
<< end >>
