magic
tech sky130A
magscale 1 2
timestamp 1702718534
<< nwell >>
rect -103 311 0 519
rect 303 311 429 519
rect 941 311 1159 519
rect 1525 311 1743 519
rect 1833 311 2051 519
rect 2452 311 2583 519
<< psubdiff >>
rect 324 75 382 99
rect 324 15 336 75
rect 370 15 382 75
rect 324 -9 382 15
<< nsubdiff >>
rect 339 445 397 469
rect 339 385 351 445
rect 385 385 397 445
rect 339 361 397 385
<< psubdiffcont >>
rect 336 15 370 75
<< nsubdiffcont >>
rect 351 385 385 445
<< poly >>
rect -52 311 8 327
rect 94 311 124 347
rect -52 277 -36 311
rect -2 277 124 311
rect -52 261 8 277
rect 94 134 124 277
rect 182 327 212 347
rect 182 311 262 327
rect 182 277 212 311
rect 246 277 262 311
rect 182 261 262 277
rect 182 134 212 261
rect 364 180 430 196
rect 511 180 541 347
rect 364 146 380 180
rect 414 146 541 180
rect 364 130 430 146
rect 511 134 541 146
rect 599 196 629 347
rect 817 335 847 347
rect 817 319 897 335
rect 817 285 847 319
rect 881 285 897 319
rect 817 269 897 285
rect 943 258 1009 274
rect 1095 258 1125 347
rect 943 224 959 258
rect 993 224 1125 258
rect 817 197 898 213
rect 943 208 1009 224
rect 599 180 679 196
rect 599 146 629 180
rect 663 146 679 180
rect 599 134 679 146
rect 817 163 847 197
rect 881 163 898 197
rect 817 146 898 163
rect 817 134 847 146
rect 1095 134 1125 224
rect 1183 325 1213 347
rect 1401 325 1431 347
rect 1709 325 1739 347
rect 1183 309 1263 325
rect 1183 275 1213 309
rect 1247 275 1263 309
rect 1183 259 1263 275
rect 1401 309 1481 325
rect 1401 275 1431 309
rect 1465 275 1481 309
rect 1401 259 1481 275
rect 1709 309 1789 325
rect 1709 275 1739 309
rect 1773 275 1789 309
rect 1709 259 1789 275
rect 1873 296 1939 312
rect 2023 296 2053 347
rect 1873 261 1889 296
rect 1923 261 2053 296
rect 1183 134 1213 259
rect 1873 245 1939 261
rect 1497 183 1563 199
rect 1497 163 1513 183
rect 1401 149 1513 163
rect 1547 149 1563 183
rect 1805 183 1871 199
rect 1805 171 1821 183
rect 613 130 679 134
rect 1401 133 1563 149
rect 1709 149 1821 171
rect 1855 149 1871 183
rect 1709 141 1871 149
rect 2023 141 2053 261
rect 2111 312 2141 347
rect 2329 335 2359 347
rect 2329 319 2409 335
rect 2111 296 2191 312
rect 2111 261 2141 296
rect 2175 261 2191 296
rect 2329 285 2359 319
rect 2393 285 2409 319
rect 2329 269 2409 285
rect 2111 245 2191 261
rect 1805 133 1871 141
rect 2111 138 2141 245
rect 2329 207 2409 223
rect 2329 173 2359 207
rect 2393 173 2409 207
rect 2329 157 2409 173
rect 2329 141 2359 157
<< polycont >>
rect -36 277 -2 311
rect 212 277 246 311
rect 380 146 414 180
rect 847 285 881 319
rect 959 224 993 258
rect 629 146 663 180
rect 847 163 881 197
rect 1213 275 1247 309
rect 1431 275 1465 309
rect 1739 275 1773 309
rect 1889 261 1923 296
rect 1513 149 1547 183
rect 1821 149 1855 183
rect 2141 261 2175 296
rect 2359 285 2393 319
rect 2359 173 2393 207
<< locali >>
rect 351 445 385 461
rect 641 399 805 433
rect 351 369 385 385
rect 893 369 993 403
rect 1225 399 1389 433
rect 1477 399 1615 433
rect 1785 399 1923 433
rect 48 311 82 369
rect -52 277 -36 311
rect -2 277 14 311
rect 48 277 212 311
rect 246 277 344 311
rect 48 112 82 277
rect 310 258 344 277
rect 465 180 499 369
rect 170 146 380 180
rect 414 146 430 180
rect 465 146 629 180
rect 663 146 679 180
rect 465 112 499 146
rect 771 112 805 369
rect 847 319 881 335
rect 847 269 881 285
rect 959 258 993 369
rect 847 197 881 213
rect 847 146 881 163
rect 959 112 993 224
rect 1049 309 1083 369
rect 1049 275 1213 309
rect 1247 275 1263 309
rect 1049 112 1083 275
rect 336 75 370 91
rect 641 50 805 84
rect 859 78 993 112
rect 1355 111 1389 369
rect 1431 309 1465 325
rect 1431 189 1465 275
rect 1513 183 1547 311
rect 1513 133 1547 149
rect 1581 258 1615 399
rect 1225 50 1389 84
rect 1581 81 1615 224
rect 1663 119 1697 369
rect 1739 309 1773 325
rect 1739 188 1773 275
rect 1821 183 1855 311
rect 1821 133 1855 149
rect 1889 296 1923 399
rect 2187 398 2283 432
rect 1889 81 1923 261
rect 1977 296 2011 374
rect 2403 369 2466 403
rect 1977 262 2141 296
rect 2011 261 2141 262
rect 2175 261 2191 296
rect 1977 119 2011 228
rect 2283 119 2317 369
rect 2359 319 2393 335
rect 2359 269 2393 285
rect 2359 207 2393 223
rect 2359 157 2393 173
rect 2432 121 2466 369
rect 2400 120 2466 121
rect 1477 47 1615 81
rect 1785 47 1923 81
rect 2187 57 2283 91
rect 2403 86 2466 120
rect 336 -1 370 15
rect 1049 -5 1083 30
rect 1663 -5 1697 27
rect 1049 -39 1697 -5
rect 1889 -5 1923 47
rect 2371 -5 2405 30
rect 1889 -39 2405 -5
<< viali >>
rect 351 398 385 432
rect -36 277 -2 311
rect 310 224 344 258
rect 136 146 170 180
rect 847 285 881 319
rect 959 224 993 258
rect 847 163 881 197
rect 336 28 370 62
rect 1431 155 1465 189
rect 1513 311 1547 345
rect 1581 224 1615 258
rect 1739 154 1773 188
rect 1821 311 1855 345
rect 1977 228 2011 262
rect 2359 285 2393 319
rect 2359 173 2393 207
<< metal1 >>
rect -103 485 2583 519
rect 136 457 170 485
rect 351 438 385 485
rect 553 457 587 485
rect 1137 445 1171 485
rect 2065 457 2099 485
rect 339 432 397 438
rect 339 398 351 432
rect 385 398 397 432
rect 339 392 397 398
rect 224 345 258 373
rect 1501 345 1559 351
rect 1809 345 1867 351
rect 224 319 1513 345
rect -48 311 10 317
rect -103 277 -36 311
rect -2 277 10 311
rect -48 271 10 277
rect 224 311 847 319
rect 124 180 182 186
rect -103 146 136 180
rect 170 146 182 180
rect 124 140 182 146
rect 224 108 258 311
rect 835 285 847 311
rect 881 311 1513 319
rect 1547 311 1821 345
rect 1855 319 2405 345
rect 1855 311 2359 319
rect 881 285 893 311
rect 1501 305 1559 311
rect 1809 305 1867 311
rect 835 279 893 285
rect 2347 285 2359 311
rect 2393 285 2405 319
rect 2347 279 2405 285
rect 298 258 356 264
rect 298 224 310 258
rect 344 224 356 258
rect 298 218 356 224
rect 947 258 1005 264
rect 1569 258 1627 264
rect 947 224 959 258
rect 993 224 1581 258
rect 1615 224 1627 258
rect 947 218 1005 224
rect 1569 218 1627 224
rect 1958 219 1968 271
rect 2020 219 2030 271
rect 2456 223 2466 275
rect 2518 266 2528 275
rect 2518 232 2583 266
rect 2518 223 2528 232
rect 310 180 344 218
rect 2346 207 2405 215
rect 835 197 893 203
rect 835 180 847 197
rect 310 163 847 180
rect 881 180 893 197
rect 1419 189 1477 195
rect 1419 180 1431 189
rect 881 163 1431 180
rect 310 155 1431 163
rect 1465 180 1477 189
rect 1727 188 1785 194
rect 1727 180 1739 188
rect 1465 155 1739 180
rect 310 154 1739 155
rect 1773 180 1785 188
rect 2346 180 2359 207
rect 1773 173 2359 180
rect 2393 173 2405 207
rect 1773 154 2405 173
rect 310 146 2405 154
rect 324 62 382 68
rect 324 28 336 62
rect 370 28 382 62
rect 136 -5 170 24
rect 324 -5 382 28
rect 553 -5 587 36
rect 1137 -5 1171 34
rect 2065 -5 2099 34
rect -103 -6 1171 -5
rect 1818 -6 2261 -5
rect -103 -39 2583 -6
<< via1 >>
rect 1968 262 2020 271
rect 1968 228 1977 262
rect 1977 228 2011 262
rect 2011 228 2020 262
rect 1968 219 2020 228
rect 2466 223 2518 275
<< metal2 >>
rect 1968 271 2020 281
rect 2466 275 2518 285
rect 2020 232 2466 266
rect 1968 209 2020 219
rect 2466 213 2518 223
use sky130_fd_pr__nfet_01v8_A6LSUL  m1
timestamp 1702713014
transform -1 0 109 0 1 66
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m2
timestamp 1702713014
transform -1 0 109 0 1 415
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_A6LSUL  m3
timestamp 1702713014
transform 1 0 197 0 1 66
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m4
timestamp 1702713014
transform 1 0 197 0 1 415
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_A6LSUL  m5
timestamp 1702713014
transform -1 0 526 0 1 66
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m6
timestamp 1702713014
transform -1 0 526 0 1 415
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m7
timestamp 1702713014
transform 1 0 614 0 1 415
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_A6LSUL  m8
timestamp 1702713014
transform 1 0 614 0 1 66
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m9
timestamp 1702713014
transform -1 0 832 0 1 415
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_A6LSUL  m10
timestamp 1702713014
transform 1 0 832 0 1 66
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m11
timestamp 1702713014
transform -1 0 1110 0 1 415
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_A6LSUL  m12
timestamp 1702713014
transform -1 0 1110 0 1 76
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m13
timestamp 1702713014
transform 1 0 1198 0 1 415
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_A6LSUL  m14
timestamp 1702713014
transform 1 0 1198 0 1 76
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m15
timestamp 1702713014
transform 1 0 1416 0 1 415
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_A6LSUL  m16
timestamp 1702713014
transform 1 0 1416 0 1 75
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m17
timestamp 1702713014
transform 1 0 1724 0 1 415
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_A6LSUL  m18
timestamp 1702713014
transform 1 0 1724 0 1 73
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m19
timestamp 1702713014
transform -1 0 2038 0 1 415
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_A6LSUL  m20
timestamp 1702713014
transform -1 0 2038 0 1 75
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m21
timestamp 1702713014
transform 1 0 2126 0 1 415
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_A6LSUL  m22
timestamp 1702713014
transform 1 0 2126 0 1 75
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m23
timestamp 1702713014
transform 1 0 2344 0 1 415
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_A6LSUL  m24
timestamp 1702713014
transform 1 0 2344 0 1 75
box -73 -68 73 68
<< labels >>
rlabel metal1 2549 232 2583 266 0 q
rlabel metal1 -103 277 -69 311 0 clk
rlabel metal1 -103 146 -69 180 0 d
rlabel metal1 -103 485 -69 519 0 VDD
rlabel metal1 -103 -39 -69 -5 0 VSS
<< end >>
