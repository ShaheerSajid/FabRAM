magic
tech sky130A
magscale 1 2
timestamp 1702289754
<< nwell >>
rect -199 60 0 268
rect 306 60 521 268
<< psubdiff >>
rect 111 -306 193 -282
rect 111 -340 136 -306
rect 170 -340 193 -306
rect 111 -364 193 -340
<< nsubdiff >>
rect 324 194 406 206
rect 324 134 348 194
rect 382 134 406 194
rect 324 122 406 134
<< psubdiffcont >>
rect 136 -340 170 -306
<< nsubdiffcont >>
rect 348 134 382 194
<< poly >>
rect 94 87 124 96
rect 58 75 124 87
rect 58 41 74 75
rect 108 41 124 75
rect 58 30 124 41
rect -172 7 -76 23
rect -172 -27 -156 7
rect -122 -27 -76 7
rect -172 -43 -76 -27
rect 94 -42 124 30
rect 182 19 212 96
rect 182 4 248 19
rect 182 -30 198 4
rect 232 -30 248 4
rect -106 -82 -76 -43
rect 182 -47 248 -30
rect 379 7 445 23
rect 379 -27 395 7
rect 429 -27 445 7
rect 379 -43 445 -27
rect 396 -82 426 -43
<< polycont >>
rect 74 41 108 75
rect -156 -27 -122 7
rect 198 -30 232 4
rect 395 -27 429 7
<< locali >>
rect 348 194 382 218
rect -10 118 82 152
rect -172 -27 -165 7
rect -113 -27 -106 7
rect -10 4 24 118
rect 224 75 258 119
rect 348 110 382 134
rect 58 41 74 75
rect 108 41 316 75
rect -64 -30 198 4
rect 232 -30 248 4
rect -64 -104 -30 -30
rect 48 -64 82 -30
rect 282 -64 316 41
rect 379 -27 386 7
rect 438 -27 445 7
rect 224 -98 384 -64
rect 350 -104 384 -98
rect 111 -306 193 -282
rect 111 -340 136 -306
rect 170 -340 193 -306
rect 111 -364 193 -340
<< viali >>
rect 348 134 382 194
rect -165 7 -113 25
rect -165 -27 -156 7
rect -156 -27 -122 7
rect -122 -27 -113 7
rect 386 7 438 25
rect 386 -27 395 7
rect 395 -27 429 7
rect 429 -27 438 7
rect 136 -340 170 -306
<< metal1 >>
rect -199 234 521 268
rect 136 206 170 234
rect 348 206 382 234
rect 342 194 388 206
rect 342 134 348 194
rect 382 134 388 194
rect 342 122 388 134
rect -177 25 -101 31
rect -177 16 -165 25
rect -199 -18 -165 16
rect -177 -27 -165 -18
rect -113 16 -101 25
rect 374 25 450 31
rect 374 16 386 25
rect -113 -18 386 16
rect -113 -27 -101 -18
rect -177 -33 -101 -27
rect 374 -27 386 -18
rect 438 16 450 25
rect 438 -18 521 16
rect 438 -27 450 -18
rect 374 -33 450 -27
rect -171 -222 -161 -170
rect -109 -222 -99 -170
rect 419 -222 429 -170
rect 481 -222 491 -170
rect 136 -256 170 -228
rect -199 -290 521 -256
rect 124 -306 183 -290
rect 124 -340 136 -306
rect 170 -340 183 -306
rect 124 -345 183 -340
rect 124 -346 182 -345
<< via1 >>
rect -161 -222 -109 -170
rect 429 -222 481 -170
<< metal2 >>
rect -161 -170 -109 300
rect -161 -381 -109 -222
rect 429 -170 481 300
rect 429 -381 481 -222
use sky130_fd_pr__pfet_01v8_4Y88KP  m1
timestamp 1702281156
transform -1 0 109 0 1 164
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m2
timestamp 1702281156
transform 1 0 197 0 1 164
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_BBXUYH  m3
timestamp 1702281156
transform -1 0 109 0 1 -148
box -73 -106 73 106
use sky130_fd_pr__nfet_01v8_BBXUYH  m4
timestamp 1702281156
transform 1 0 197 0 1 -148
box -73 -106 73 106
use sky130_fd_pr__nfet_01v8_FB3UY2  m5
timestamp 1702281156
transform 1 0 -91 0 1 -168
box -73 -86 73 86
use sky130_fd_pr__nfet_01v8_FB3UY2  m6
timestamp 1702281156
transform 1 0 411 0 1 -168
box -73 -86 73 86
<< labels >>
rlabel metal2 -161 268 -109 300 1 BL
rlabel metal1 -199 234 -161 268 1 VDD
rlabel metal1 -199 -18 -177 16 1 WL
rlabel metal1 -199 -290 -161 -256 1 VSS
rlabel metal2 429 268 481 300 1 BL_
<< end >>
