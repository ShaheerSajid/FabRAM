magic
tech sky130A
magscale 1 2
timestamp 1702461067
<< metal1 >>
rect 0 262 196 296
rect 161 -291 196 262
rect 637 -91 647 -39
rect 699 -91 709 -39
rect 969 -285 979 -282
rect 161 -325 685 -291
rect 967 -331 979 -285
rect 969 -334 979 -331
rect 1031 -334 1041 -282
rect 1299 -285 1309 -282
rect 1297 -331 1309 -285
rect 1299 -334 1309 -331
rect 1361 -334 1371 -282
rect 557 -597 567 -545
rect 619 -563 629 -545
rect 619 -597 685 -563
<< via1 >>
rect 647 -91 699 -39
rect 979 -334 1031 -282
rect 1309 -334 1361 -282
rect 567 -597 619 -545
<< metal2 >>
rect 567 -545 619 0
rect 567 -674 619 -597
rect 647 -39 699 0
rect 647 -674 699 -91
rect 977 -280 1033 -270
rect 977 -346 1033 -336
rect 1307 -280 1363 -270
rect 1307 -346 1363 -336
<< via2 >>
rect 977 -282 1033 -280
rect 977 -334 979 -282
rect 979 -334 1031 -282
rect 1031 -334 1033 -282
rect 977 -336 1033 -334
rect 1307 -282 1363 -280
rect 1307 -334 1309 -282
rect 1309 -334 1361 -282
rect 1361 -334 1363 -282
rect 1307 -336 1363 -334
<< metal3 >>
rect 967 -280 1132 -275
rect 967 -336 977 -280
rect 1033 -336 1132 -280
rect 967 -341 1132 -336
rect 1297 -280 1462 -275
rect 1297 -336 1307 -280
rect 1363 -336 1462 -280
rect 1297 -341 1462 -336
rect 1066 -652 1132 -341
rect 1066 -718 1462 -652
use dec_2to4  dec_2to4_0 ~/Desktop/FabRAM/FE/sram130/dec_2to4
timestamp 1702458901
transform 1 0 0 0 1 0
box 0 0 1462 2422
use not  not_0 ~/Desktop/FabRAM/FE/sram130/not
timestamp 1702458901
transform 1 0 685 0 1 -688
box 0 91 330 649
use not  not_1
timestamp 1702458901
transform 1 0 1015 0 1 -688
box 0 91 330 649
<< labels >>
rlabel via1 1311 -325 1345 -291 0 B
rlabel via1 981 -325 1015 -291 0 B
rlabel metal3 1066 -341 1132 -275 0 Y3
rlabel metal3 1396 -341 1462 -275 0 Y3
<< end >>
