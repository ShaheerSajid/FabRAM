magic
tech sky130A
magscale 1 2
timestamp 1702386201
<< poly >>
rect 94 472 124 477
rect 44 456 124 472
rect 44 422 60 456
rect 94 422 124 456
rect 44 406 124 422
rect 94 264 124 406
rect 182 401 212 477
rect 170 385 224 401
rect 170 351 180 385
rect 214 351 224 385
rect 170 335 224 351
rect 182 264 212 335
rect 270 326 300 477
rect 270 310 350 326
rect 270 276 300 310
rect 334 276 350 310
rect 270 264 350 276
rect 300 260 350 264
<< polycont >>
rect 60 422 94 456
rect 180 351 214 385
rect 300 276 334 310
<< locali >>
rect 44 422 60 456
rect 94 422 110 456
rect 164 351 180 385
rect 214 351 230 385
rect 164 276 180 310
rect 214 276 300 310
rect 334 276 350 310
<< viali >>
rect 60 422 94 456
rect 180 351 214 385
rect 180 276 214 310
<< metal1 >>
rect 0 615 394 649
rect 48 587 82 615
rect 224 587 258 615
rect 136 475 170 503
rect 312 475 346 503
rect 48 456 106 462
rect 0 422 60 456
rect 94 422 106 456
rect 136 441 346 475
rect 48 416 106 422
rect 312 397 346 441
rect 168 385 226 391
rect 0 351 180 385
rect 214 351 226 385
rect 168 345 226 351
rect 312 363 394 397
rect 168 310 226 316
rect 0 276 180 310
rect 214 276 226 310
rect 168 270 226 276
rect 312 238 346 363
rect 48 125 82 154
rect 0 91 394 125
use sky130_fd_pr__nfet_01v8_A6LSUL  m1 ~/Desktop/FabRAM/FE/sram130/common
timestamp 1702353901
transform 1 0 109 0 1 196
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_A6LSUL  m2
timestamp 1702353901
transform 1 0 197 0 1 196
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_A6LSUL  m3
timestamp 1702353901
transform 1 0 285 0 1 196
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m4 ~/Desktop/FabRAM/FE/sram130/common
timestamp 1702353901
transform 1 0 109 0 1 545
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m5
timestamp 1702353901
transform -1 0 197 0 1 545
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m6
timestamp 1702353901
transform 1 0 285 0 1 545
box -109 -104 109 104
<< labels >>
rlabel metal1 0 615 34 649 0 VDD
rlabel metal1 0 422 34 456 0 A
rlabel metal1 0 351 34 385 0 B
rlabel metal1 0 276 34 310 0 C
rlabel metal1 0 91 34 125 0 VSS
rlabel metal1 360 363 394 397 0 Y
<< end >>
