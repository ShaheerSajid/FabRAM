magic
tech sky130A
magscale 1 2
timestamp 1703829263
<< metal1 >>
rect 154 2173 164 2195
rect 0 2139 164 2173
rect 220 2139 230 2195
rect 248 1477 258 1499
rect 0 1443 258 1477
rect 314 1443 324 1499
rect 1348 1042 1382 2425
rect 1348 1008 1458 1042
rect 332 781 342 803
rect 0 747 342 781
rect 398 747 408 803
rect 426 85 436 107
rect 0 51 436 85
rect 492 51 502 107
<< via1 >>
rect 164 2139 220 2195
rect 258 1443 314 1499
rect 342 747 398 803
rect 436 51 492 107
<< metal2 >>
rect 164 2295 220 2305
rect 164 2195 220 2239
rect 164 2088 220 2139
rect 258 2169 314 2179
rect 258 1499 314 2113
rect 258 1392 314 1443
rect 342 2043 398 2053
rect 342 803 398 1987
rect 342 696 398 747
rect 436 1917 492 1927
rect 436 107 492 1861
rect 436 0 492 51
<< via2 >>
rect 164 2239 220 2295
rect 258 2113 314 2169
rect 342 1987 398 2043
rect 436 1861 492 1917
<< metal3 >>
rect 154 2295 1458 2300
rect 154 2239 164 2295
rect 220 2239 1458 2295
rect 154 2234 1458 2239
rect 248 2169 1458 2174
rect 248 2113 258 2169
rect 314 2113 1458 2169
rect 248 2108 1458 2113
rect 332 2043 1458 2048
rect 332 1987 342 2043
rect 398 1987 1458 2043
rect 332 1982 1458 1987
rect 426 1917 1458 1922
rect 426 1861 436 1917
rect 492 1861 1458 1917
rect 426 1856 1458 1861
<< end >>
