magic
tech sky130A
magscale 1 2
timestamp 1702726551
<< nwell >>
rect 306 -338 339 -130
rect 0 -425 339 -338
rect 643 -425 720 -130
rect 187 -1412 327 -1088
<< psubdiff >>
rect 237 580 319 604
rect 237 546 262 580
rect 296 546 319 580
rect 237 522 319 546
<< nsubdiff >>
rect 223 -1226 305 -1214
rect 223 -1286 247 -1226
rect 281 -1286 305 -1226
rect 223 -1298 305 -1286
<< psubdiffcont >>
rect 262 546 296 580
<< nsubdiffcont >>
rect 247 -1286 281 -1226
<< poly >>
rect 94 556 193 572
rect 94 522 143 556
rect 177 522 193 556
rect 94 506 193 522
rect 94 479 125 506
rect 262 247 328 258
rect 262 233 278 247
rect 182 213 278 233
rect 312 213 328 247
rect 182 203 328 213
rect 39 160 124 176
rect 39 126 55 160
rect 89 126 124 160
rect 39 110 124 126
rect 94 49 124 110
rect 182 49 212 203
rect 286 133 352 149
rect 432 133 462 179
rect 286 99 302 133
rect 336 99 462 133
rect 286 83 352 99
rect 432 63 462 99
rect 520 174 550 179
rect 520 158 600 174
rect 520 124 550 158
rect 584 124 600 158
rect 520 109 600 124
rect 520 63 550 109
rect 94 -338 212 -302
rect 120 -372 136 -338
rect 170 -372 186 -338
rect 120 -388 186 -372
rect 421 -1397 451 -1376
rect 538 -1397 593 -1381
rect 421 -1431 549 -1397
rect 583 -1431 593 -1397
rect 421 -1454 451 -1431
rect 538 -1447 593 -1431
<< polycont >>
rect 143 522 177 556
rect 278 213 312 247
rect 55 126 89 160
rect 302 99 336 133
rect 550 124 584 158
rect 136 -372 170 -338
rect 549 -1431 583 -1397
<< locali >>
rect 143 556 177 739
rect 237 580 319 604
rect 237 546 262 580
rect 296 546 319 580
rect 237 522 319 546
rect 143 506 177 522
rect 262 213 278 247
rect 312 213 328 247
rect 562 201 668 235
rect 39 126 55 160
rect 89 126 105 160
rect 386 158 420 201
rect 224 99 302 133
rect 336 99 352 133
rect 386 124 550 158
rect 584 124 600 158
rect 224 27 258 99
rect 386 41 420 124
rect 634 42 668 201
rect 562 8 668 42
rect 48 -188 82 -65
rect 224 -188 258 -65
rect 48 -338 82 -280
rect 48 -372 136 -338
rect 170 -372 186 -338
rect 386 -411 420 -367
rect 46 -445 420 -411
rect 46 -522 80 -445
rect 247 -1226 281 -1202
rect 281 -1272 375 -1238
rect 247 -1310 281 -1286
rect 549 -1397 583 -925
rect 549 -1452 583 -1431
<< viali >>
rect 143 739 177 773
rect 262 546 296 580
rect 278 213 312 247
rect 55 126 89 160
rect 46 -556 80 -522
<< metal1 >>
rect 316 865 326 883
rect 12 831 326 865
rect 378 865 388 883
rect 378 831 720 865
rect 131 773 189 779
rect 234 773 244 791
rect 12 739 143 773
rect 177 739 244 773
rect 296 773 306 791
rect 296 739 720 773
rect 131 733 189 739
rect 396 678 406 696
rect 12 644 406 678
rect 458 678 468 696
rect 458 644 720 678
rect 48 453 82 644
rect 237 580 309 644
rect 474 605 508 644
rect 237 546 262 580
rect 296 546 309 580
rect 237 522 309 546
rect 36 117 46 169
rect 98 117 108 169
rect 136 23 170 285
rect 266 247 324 253
rect 266 213 278 247
rect 312 213 324 247
rect 266 207 324 213
rect 278 152 312 207
rect 630 152 640 161
rect 278 118 640 152
rect 630 109 640 118
rect 692 109 702 161
rect 135 -459 170 -276
rect 380 -363 390 -310
rect 602 -362 628 -310
rect 680 -362 690 -310
rect 602 -363 690 -362
rect 316 -459 326 -407
rect 378 -459 388 -407
rect 474 -459 509 -363
rect 27 -565 37 -513
rect 90 -565 100 -513
rect 234 -711 244 -659
rect 296 -711 306 -659
rect 396 -983 406 -949
rect 249 -1480 283 -983
rect 382 -1001 406 -983
rect 458 -1001 468 -949
rect 316 -1133 326 -1080
rect 378 -1133 415 -1080
rect 316 -1150 415 -1133
rect 463 -1480 497 -1338
rect 249 -1514 409 -1480
rect 463 -1749 497 -1680
<< via1 >>
rect 326 831 378 883
rect 244 739 296 791
rect 406 644 458 696
rect 46 160 98 169
rect 46 126 55 160
rect 55 126 89 160
rect 89 126 98 160
rect 46 117 98 126
rect 640 109 692 161
rect 628 -362 680 -310
rect 326 -459 378 -407
rect 37 -522 90 -513
rect 37 -556 46 -522
rect 46 -556 80 -522
rect 80 -556 90 -522
rect 37 -565 90 -556
rect 244 -711 296 -659
rect 406 -1001 458 -949
rect 326 -1133 378 -1080
<< metal2 >>
rect 12 719 64 917
rect 12 685 98 719
rect 46 169 98 685
rect 46 107 98 117
rect 37 -513 90 -503
rect 37 -575 90 -565
rect 164 -1749 216 917
rect 326 883 378 890
rect 244 791 296 801
rect 244 -659 296 739
rect 244 -721 296 -711
rect 326 -407 378 831
rect 326 -1080 378 -459
rect 406 696 458 706
rect 406 -949 458 644
rect 406 -1011 458 -1001
rect 326 -1143 378 -1133
rect 488 -1749 540 918
rect 640 161 692 917
rect 640 99 692 109
rect 628 -310 680 -300
rect 628 -425 680 -362
use bit_cell  bit_cell_0 ~/Desktop/FabRAM/FE/sram130/bit_cell
timestamp 1702653557
transform 1 0 0 0 1 -1121
box 0 0 720 696
use sky130_fd_pr__nfet_01v8_A6LSUL  m1
timestamp 1702653557
transform -1 0 109 0 1 -19
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_A6LSUL  m2
timestamp 1702653557
transform 1 0 197 0 1 -19
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP#0  m3
timestamp 1702552054
transform -1 0 109 0 1 -234
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP#0  m4
timestamp 1702552054
transform 1 0 197 0 1 -234
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_5YUHNA  m5
timestamp 1702553317
transform -1 0 447 0 1 -163
box -109 -262 109 262
use sky130_fd_pr__nfet_01v8_JB3UY8  m6
timestamp 1702553317
transform -1 0 447 0 1 405
box -73 -226 73 226
use sky130_fd_pr__pfet_01v8_5YUHNA  m7
timestamp 1702553317
transform 1 0 535 0 1 -163
box -109 -262 109 262
use sky130_fd_pr__nfet_01v8_JB3UY8  m8
timestamp 1702553317
transform 1 0 535 0 1 405
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_VJ5ZNR  m9
timestamp 1702559342
transform 1 0 109 0 1 369
box -73 -110 73 110
use sky130_fd_pr__nfet_01v8_L8ATA9  m10
timestamp 1702726551
transform 1 0 436 0 1 -1580
box -73 -126 73 126
use sky130_fd_pr__pfet_01v8_5SMHNA  m11
timestamp 1702726551
transform 1 0 436 0 1 -1250
box -109 -162 109 162
<< labels >>
rlabel metal2 12 865 64 917 0 DR_
rlabel metal2 164 865 216 917 0 DW_
rlabel metal2 488 866 540 918 0 DW
rlabel metal2 640 865 692 917 0 DR
rlabel metal1 12 831 46 865 0 VDD
rlabel metal1 12 739 46 773 0 SAEN
rlabel metal1 12 644 46 678 0 VSS
rlabel space 0 -459 34 -425 0 VDD
rlabel space 0 -983 34 -949 0 VSS
rlabel metal2 164 -1749 216 -1697 0 DW_
rlabel metal2 488 -1749 540 -1697 0 DW
rlabel metal1 463 -1749 497 -1715 0 SB
<< end >>
