magic
tech sky130A
magscale 1 2
timestamp 1702452662
<< nwell >>
rect 0 488 876 696
<< nmos >>
rect 94 201 124 285
rect 182 201 212 285
rect 400 201 430 285
rect 488 201 518 285
rect 576 201 606 285
rect 664 201 694 285
rect 752 201 782 285
<< pmos >>
rect 94 550 124 634
rect 182 550 212 634
rect 400 550 430 634
rect 488 550 518 634
rect 576 550 606 634
rect 664 550 694 634
rect 752 550 782 634
<< ndiff >>
rect 36 273 94 285
rect 36 213 48 273
rect 82 213 94 273
rect 36 201 94 213
rect 124 273 182 285
rect 124 213 136 273
rect 170 213 182 273
rect 124 201 182 213
rect 212 273 270 285
rect 212 213 224 273
rect 258 213 270 273
rect 212 201 270 213
rect 342 273 400 285
rect 342 213 354 273
rect 388 213 400 273
rect 342 201 400 213
rect 430 273 488 285
rect 430 213 442 273
rect 476 213 488 273
rect 430 201 488 213
rect 518 273 576 285
rect 518 213 530 273
rect 564 213 576 273
rect 518 201 576 213
rect 606 273 664 285
rect 606 213 618 273
rect 652 213 664 273
rect 606 201 664 213
rect 694 273 752 285
rect 694 213 706 273
rect 740 213 752 273
rect 694 201 752 213
rect 782 273 840 285
rect 782 213 794 273
rect 828 213 840 273
rect 782 201 840 213
<< pdiff >>
rect 36 622 94 634
rect 36 562 48 622
rect 82 562 94 622
rect 36 550 94 562
rect 124 622 182 634
rect 124 562 136 622
rect 170 562 182 622
rect 124 550 182 562
rect 212 622 270 634
rect 212 562 224 622
rect 258 562 270 622
rect 212 550 270 562
rect 342 622 400 634
rect 342 562 354 622
rect 388 562 400 622
rect 342 550 400 562
rect 430 622 488 634
rect 430 562 442 622
rect 476 562 488 622
rect 430 550 488 562
rect 518 622 576 634
rect 518 562 530 622
rect 564 562 576 622
rect 518 550 576 562
rect 606 622 664 634
rect 606 562 618 622
rect 652 562 664 622
rect 606 550 664 562
rect 694 622 752 634
rect 694 562 706 622
rect 740 562 752 622
rect 694 550 752 562
rect 782 622 840 634
rect 782 562 794 622
rect 828 562 840 622
rect 782 550 840 562
<< ndiffc >>
rect 48 213 82 273
rect 136 213 170 273
rect 224 213 258 273
rect 354 213 388 273
rect 442 213 476 273
rect 530 213 564 273
rect 618 213 652 273
rect 706 213 740 273
rect 794 213 828 273
<< pdiffc >>
rect 48 562 82 622
rect 136 562 170 622
rect 224 562 258 622
rect 354 562 388 622
rect 442 562 476 622
rect 530 562 564 622
rect 618 562 652 622
rect 706 562 740 622
rect 794 562 828 622
<< poly >>
rect 94 634 124 660
rect 182 634 212 660
rect 400 634 430 660
rect 488 634 518 660
rect 576 634 606 660
rect 664 634 694 660
rect 752 634 782 660
rect 94 518 124 550
rect 44 502 124 518
rect 44 468 60 502
rect 94 468 124 502
rect 44 452 124 468
rect 94 285 124 452
rect 182 373 212 550
rect 400 462 430 550
rect 347 444 430 462
rect 488 444 518 550
rect 576 444 606 550
rect 664 444 694 550
rect 752 444 782 550
rect 347 410 357 444
rect 391 410 782 444
rect 347 394 430 410
rect 182 357 262 373
rect 182 323 212 357
rect 246 323 262 357
rect 182 307 262 323
rect 182 285 212 307
rect 400 285 430 394
rect 488 285 518 410
rect 576 285 606 410
rect 664 285 694 410
rect 752 285 782 410
rect 94 175 124 201
rect 182 175 212 201
rect 400 175 430 201
rect 488 175 518 201
rect 576 175 606 201
rect 664 175 694 201
rect 752 175 782 201
<< polycont >>
rect 60 468 94 502
rect 357 410 391 444
rect 212 323 246 357
<< locali >>
rect 48 622 82 638
rect 48 546 82 562
rect 136 622 170 638
rect 136 546 170 562
rect 224 622 258 638
rect 224 546 258 562
rect 354 622 388 638
rect 354 546 388 562
rect 442 622 476 638
rect 44 468 60 502
rect 94 468 110 502
rect 442 496 476 562
rect 530 622 564 638
rect 530 546 564 562
rect 618 622 652 638
rect 618 496 652 562
rect 706 622 740 638
rect 706 546 740 562
rect 794 622 828 638
rect 794 496 828 562
rect 442 461 828 496
rect 794 444 828 461
rect 340 410 357 444
rect 391 410 407 444
rect 794 358 828 410
rect 48 323 60 357
rect 94 323 212 357
rect 246 323 262 357
rect 442 323 828 358
rect 48 273 82 289
rect 48 197 82 213
rect 136 273 170 289
rect 136 197 170 213
rect 224 273 258 289
rect 224 197 258 213
rect 354 273 388 289
rect 354 197 388 213
rect 442 273 476 323
rect 442 197 476 213
rect 530 273 564 289
rect 530 197 564 213
rect 618 273 652 323
rect 618 197 652 213
rect 706 273 740 289
rect 706 197 740 213
rect 794 273 828 323
rect 794 197 828 213
<< viali >>
rect 48 562 82 622
rect 136 562 170 622
rect 224 562 258 622
rect 354 562 388 622
rect 442 562 476 622
rect 60 468 94 502
rect 530 562 564 622
rect 618 562 652 622
rect 706 562 740 622
rect 794 562 828 622
rect 357 410 391 444
rect 794 410 828 444
rect 60 323 94 357
rect 48 213 82 273
rect 136 213 170 273
rect 224 213 258 273
rect 354 213 388 273
rect 442 213 476 273
rect 530 213 564 273
rect 618 213 652 273
rect 706 213 740 273
rect 794 213 828 273
<< metal1 >>
rect 0 662 876 696
rect 48 634 82 662
rect 224 634 258 662
rect 354 634 388 662
rect 530 634 564 662
rect 706 634 740 662
rect 42 622 88 634
rect 42 562 48 622
rect 82 562 88 622
rect 42 550 88 562
rect 130 622 176 634
rect 130 562 136 622
rect 170 562 176 622
rect 130 550 176 562
rect 218 622 264 634
rect 218 562 224 622
rect 258 562 264 622
rect 218 550 264 562
rect 348 622 394 634
rect 348 562 354 622
rect 388 562 394 622
rect 348 550 394 562
rect 436 622 482 634
rect 436 562 442 622
rect 476 562 482 622
rect 436 550 482 562
rect 524 622 570 634
rect 524 562 530 622
rect 564 562 570 622
rect 524 550 570 562
rect 612 622 658 634
rect 612 562 618 622
rect 652 562 658 622
rect 612 550 658 562
rect 700 622 746 634
rect 700 562 706 622
rect 740 562 746 622
rect 700 550 746 562
rect 788 622 834 634
rect 788 562 794 622
rect 828 562 834 622
rect 788 550 834 562
rect 48 502 106 508
rect 0 468 60 502
rect 94 468 106 502
rect 0 462 106 468
rect 0 410 34 462
rect 136 444 170 550
rect 345 444 403 450
rect 136 410 357 444
rect 391 410 403 444
rect 35 314 45 366
rect 97 314 107 366
rect 136 285 170 410
rect 345 404 403 410
rect 782 444 840 450
rect 782 410 794 444
rect 828 410 876 444
rect 782 404 840 410
rect 42 273 88 285
rect 42 213 48 273
rect 82 213 88 273
rect 42 201 88 213
rect 130 273 176 285
rect 130 213 136 273
rect 170 213 176 273
rect 130 201 176 213
rect 218 273 264 285
rect 218 213 224 273
rect 258 213 264 273
rect 218 201 264 213
rect 348 273 394 285
rect 348 213 354 273
rect 388 213 394 273
rect 348 201 394 213
rect 436 273 482 285
rect 436 213 442 273
rect 476 213 482 273
rect 436 201 482 213
rect 524 273 570 285
rect 524 213 530 273
rect 564 213 570 273
rect 524 201 570 213
rect 612 273 658 285
rect 612 213 618 273
rect 652 213 658 273
rect 612 201 658 213
rect 700 273 746 285
rect 700 213 706 273
rect 740 213 746 273
rect 700 201 746 213
rect 788 273 834 285
rect 788 213 794 273
rect 828 213 834 273
rect 788 201 834 213
rect 48 172 82 201
rect 224 172 258 201
rect 354 172 388 201
rect 530 172 564 201
rect 706 172 740 201
rect 0 138 876 172
<< via1 >>
rect 45 357 97 366
rect 45 323 60 357
rect 60 323 94 357
rect 94 323 97 357
rect 45 314 97 323
<< metal2 >>
rect 45 366 97 696
rect 45 0 97 314
<< labels >>
rlabel metal1 0 662 34 696 0 VDD
rlabel metal1 0 410 34 444 0 A
rlabel metal1 0 138 34 172 0 VSS
rlabel metal2 45 0 97 52 0 WLEN
rlabel metal1 842 410 876 444 0 B
<< end >>
