magic
tech sky130A
magscale 1 2
timestamp 1703829772
<< metal1 >>
rect 154 4957 164 4979
rect 0 4923 164 4957
rect 220 4923 230 4979
rect 248 4261 258 4283
rect 0 4227 258 4261
rect 314 4227 324 4283
rect 332 3565 342 3587
rect 0 3531 342 3565
rect 398 3531 408 3587
rect 1348 3323 1382 5209
rect 1348 3289 1458 3323
rect 426 2869 436 2891
rect 0 2835 436 2869
rect 492 2835 502 2891
rect 510 2173 520 2195
rect 0 2139 520 2173
rect 576 2139 586 2195
rect 0 1443 672 1477
rect 713 781 723 803
rect 0 747 723 781
rect 779 747 789 803
rect 811 85 821 107
rect 0 51 821 85
rect 877 51 887 107
<< via1 >>
rect 164 4923 220 4979
rect 258 4227 314 4283
rect 342 3531 398 3587
rect 436 2835 492 2891
rect 520 2139 576 2195
rect 723 747 779 803
rect 821 51 877 107
<< metal2 >>
rect 164 5079 220 5089
rect 164 4979 220 5023
rect 164 4872 220 4923
rect 258 4953 314 4963
rect 258 4283 314 4897
rect 258 4176 314 4227
rect 342 4827 398 4837
rect 342 3587 398 4771
rect 342 3480 398 3531
rect 436 4701 492 4711
rect 436 2891 492 4645
rect 436 2784 492 2835
rect 520 4575 576 4585
rect 520 4509 576 4519
rect 520 2205 575 4509
rect 616 4449 672 4459
rect 520 2195 576 2205
rect 520 2129 576 2139
rect 520 2098 575 2129
rect 616 1392 672 4393
rect 723 4323 779 4333
rect 723 803 779 4267
rect 723 696 779 747
rect 821 4197 877 4207
rect 821 107 877 4141
rect 821 0 877 51
<< via2 >>
rect 164 5023 220 5079
rect 258 4897 314 4953
rect 342 4771 398 4827
rect 436 4645 492 4701
rect 520 4519 576 4575
rect 616 4393 672 4449
rect 723 4267 779 4323
rect 821 4141 877 4197
<< metal3 >>
rect 154 5079 1458 5084
rect 154 5023 164 5079
rect 220 5023 1458 5079
rect 154 5018 1458 5023
rect 248 4953 1458 4958
rect 248 4897 258 4953
rect 314 4897 1458 4953
rect 248 4892 1458 4897
rect 332 4827 1458 4832
rect 332 4771 342 4827
rect 398 4771 1458 4827
rect 332 4766 1458 4771
rect 426 4701 1458 4706
rect 426 4645 436 4701
rect 492 4645 1458 4701
rect 426 4640 1458 4645
rect 510 4575 1458 4580
rect 510 4519 520 4575
rect 576 4519 1458 4575
rect 510 4514 1458 4519
rect 606 4449 1458 4454
rect 606 4393 616 4449
rect 672 4393 1458 4449
rect 606 4388 1458 4393
rect 713 4323 1458 4328
rect 713 4267 723 4323
rect 779 4267 1458 4323
rect 713 4262 1458 4267
rect 811 4197 1458 4202
rect 811 4141 821 4197
rect 877 4141 1458 4197
rect 811 4136 1458 4141
<< end >>
