.title sram_gen
.subckt bit_cell VDD VSS WL BL BL_
X0 Q Q_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X1 Q_ Q VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X2 Q Q_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 Q_ Q VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 Q WL BL VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
X5 Q_ WL BL_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
.ends bit_cell

.subckt dmy_cell VDD VSS WL BL BL_
X0 Q VSS VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X1 Q_ VDD VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X2 Q VSS VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 Q_ VDD VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 Q WL BL VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
X5 Q_ WL BL_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
.ends dmy_cell

.subckt in_reg VDD VSS clk D Q
X0 net3 clk VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X8 net3 clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 net4 net2 net5 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X10 Din net2 net1 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 net55 Q VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X13 net55 Q VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 net2 net3 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X11 net2 net3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X5 Din net3 net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X15 net4 net3 net5 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 Q net5 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X9 Q net5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X6 net11 net4 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X12 net11 net4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X7 net4 net1 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X14 net4 net1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X16 net11 net2 net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X17 net11 net3 net1 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X18 net55 net3 net5 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X19 net55 net2 net5 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X20 D_ D VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X21 D_ D VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X22 Din D_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X23 Din D_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
.ends in_reg

.subckt se_cell VDD VSS SAEN BL BL_ SB
X0 net1 SAEN VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.84
X1 diff1 BL_ net1 net1 sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X2 diff2 BL net1 net1 sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X3 diff1 diff1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 diff2 diff1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X5 diff2_ diff2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X6 diff2_ diff2 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=2
X7 SB_ diff2_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X8 SB_ diff2_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=2
X9 SB_w Q_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X10 Q_ SB_w VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X11 SB_w Q_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X12 Q_ SB_w VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X13 SB_w SAEN SB_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
X14 Q_ SAEN diff2_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
X15 SB SB_w VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X16 SB SB_w VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
.ends se_cell

.subckt not VDD VSS A B
X0 B A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 B A VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends not

.subckt notdel VDD VSS A B
X0 B A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.84
X1 B A VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends notdel

.subckt nand2 VDD VSS A B Y
X0 Y A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 Y B VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 Y B net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X3 net1 A VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends nand2

.subckt nand3 VDD VSS A B C Y
X0 Y A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 Y B VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 Y C VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 Y A net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X4 net1 B net2 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X5 net2 C VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends nand3

.subckt nand4 VDD VSS A B C D Y
X0 Y A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 Y B VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 Y C VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 Y D VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 Y D net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X5 net1 B net2 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X6 net2 C net3 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X7 net3 A VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends nand4

.subckt dec_2to4 VDD VSS A1 A0 Y0 Y1 Y2 Y3
X0 VDD VSS A1 A_1 not
X1 VDD VSS A0 A_0 not
X2 VDD VSS A_1 A_0 Y0_ nand2
X3 VDD VSS A_1 A0 Y1_ nand2
X4 VDD VSS A1 A_0 Y2_ nand2
X5 VDD VSS A1 A0 Y3_ nand2
X6 VDD VSS Y0_ Y0 not
X7 VDD VSS Y1_ Y1 not
X8 VDD VSS Y2_ Y2 not
X9 VDD VSS Y3_ Y3 not
.ends dec_2to4

.subckt dec_3to6 VDD VSS A2 A1 A0 Y0 Y1 Y2 Y3 Y4 Y5
X0 VDD VSS A2 Y4 not
X1 VDD VSS Y4 Y5 not
X2 VDD VSS A1 A0 Y0 Y1 Y2 Y3 dec_2to4
.ends dec_3to6

.subckt row_dec64 VDD VSS A0 A1 A2 A3 A4 A5 DC0 DC1 DC2 DC3 DC4 DC5 DC6 DC7 DC8 DC9 DC10 DC11 DC12 DC13 DC14 DC15 DC16 DC17 DC18 DC19 DC20 DC21 DC22 DC23 DC24 DC25 DC26 DC27 DC28 DC29 DC30 DC31 DC32 DC33 DC34 DC35 DC36 DC37 DC38 DC39 DC40 DC41 DC42 DC43 DC44 DC45 DC46 DC47 DC48 DC49 DC50 DC51 DC52 DC53 DC54 DC55 DC56 DC57 DC58 DC59 DC60 DC61 DC62 DC63
X0 VDD VSS A1 A0 Y0 Y1 Y2 Y3 dec_2to4
X1 VDD VSS A3 A2 Y4 Y5 Y6 Y7 dec_2to4
X2 VDD VSS A5 A4 Y8 Y9 Y10 Y11 dec_2to4
X3 VDD VSS Y0 Y4 Y8 DC_0 nand3
X4 VDD VSS Y1 Y4 Y8 DC_1 nand3
X5 VDD VSS Y2 Y4 Y8 DC_2 nand3
X6 VDD VSS Y3 Y4 Y8 DC_3 nand3
X7 VDD VSS Y0 Y5 Y8 DC_4 nand3
X8 VDD VSS Y1 Y5 Y8 DC_5 nand3
X9 VDD VSS Y2 Y5 Y8 DC_6 nand3
X10 VDD VSS Y3 Y5 Y8 DC_7 nand3
X11 VDD VSS Y0 Y6 Y8 DC_8 nand3
X12 VDD VSS Y1 Y6 Y8 DC_9 nand3
X13 VDD VSS Y2 Y6 Y8 DC_10 nand3
X14 VDD VSS Y3 Y6 Y8 DC_11 nand3
X15 VDD VSS Y0 Y7 Y8 DC_12 nand3
X16 VDD VSS Y1 Y7 Y8 DC_13 nand3
X17 VDD VSS Y2 Y7 Y8 DC_14 nand3
X18 VDD VSS Y3 Y7 Y8 DC_15 nand3
X19 VDD VSS Y0 Y4 Y9 DC_16 nand3
X20 VDD VSS Y1 Y4 Y9 DC_17 nand3
X21 VDD VSS Y2 Y4 Y9 DC_18 nand3
X22 VDD VSS Y3 Y4 Y9 DC_19 nand3
X23 VDD VSS Y0 Y5 Y9 DC_20 nand3
X24 VDD VSS Y1 Y5 Y9 DC_21 nand3
X25 VDD VSS Y2 Y5 Y9 DC_22 nand3
X26 VDD VSS Y3 Y5 Y9 DC_23 nand3
X27 VDD VSS Y0 Y6 Y9 DC_24 nand3
X28 VDD VSS Y1 Y6 Y9 DC_25 nand3
X29 VDD VSS Y2 Y6 Y9 DC_26 nand3
X30 VDD VSS Y3 Y6 Y9 DC_27 nand3
X31 VDD VSS Y0 Y7 Y9 DC_28 nand3
X32 VDD VSS Y1 Y7 Y9 DC_29 nand3
X33 VDD VSS Y2 Y7 Y9 DC_30 nand3
X34 VDD VSS Y3 Y7 Y9 DC_31 nand3
X35 VDD VSS Y0 Y4 Y10 DC_32 nand3
X36 VDD VSS Y1 Y4 Y10 DC_33 nand3
X37 VDD VSS Y2 Y4 Y10 DC_34 nand3
X38 VDD VSS Y3 Y4 Y10 DC_35 nand3
X39 VDD VSS Y0 Y5 Y10 DC_36 nand3
X40 VDD VSS Y1 Y5 Y10 DC_37 nand3
X41 VDD VSS Y2 Y5 Y10 DC_38 nand3
X42 VDD VSS Y3 Y5 Y10 DC_39 nand3
X43 VDD VSS Y0 Y6 Y10 DC_40 nand3
X44 VDD VSS Y1 Y6 Y10 DC_41 nand3
X45 VDD VSS Y2 Y6 Y10 DC_42 nand3
X46 VDD VSS Y3 Y6 Y10 DC_43 nand3
X47 VDD VSS Y0 Y7 Y10 DC_44 nand3
X48 VDD VSS Y1 Y7 Y10 DC_45 nand3
X49 VDD VSS Y2 Y7 Y10 DC_46 nand3
X50 VDD VSS Y3 Y7 Y10 DC_47 nand3
X51 VDD VSS Y0 Y4 Y11 DC_48 nand3
X52 VDD VSS Y1 Y4 Y11 DC_49 nand3
X53 VDD VSS Y2 Y4 Y11 DC_50 nand3
X54 VDD VSS Y3 Y4 Y11 DC_51 nand3
X55 VDD VSS Y0 Y5 Y11 DC_52 nand3
X56 VDD VSS Y1 Y5 Y11 DC_53 nand3
X57 VDD VSS Y2 Y5 Y11 DC_54 nand3
X58 VDD VSS Y3 Y5 Y11 DC_55 nand3
X59 VDD VSS Y0 Y6 Y11 DC_56 nand3
X60 VDD VSS Y1 Y6 Y11 DC_57 nand3
X61 VDD VSS Y2 Y6 Y11 DC_58 nand3
X62 VDD VSS Y3 Y6 Y11 DC_59 nand3
X63 VDD VSS Y0 Y7 Y11 DC_60 nand3
X64 VDD VSS Y1 Y7 Y11 DC_61 nand3
X65 VDD VSS Y2 Y7 Y11 DC_62 nand3
X66 VDD VSS Y3 Y7 Y11 DC_63 nand3
X67 VDD VSS DC_0 DC0 not
X68 VDD VSS DC_1 DC1 not
X69 VDD VSS DC_2 DC2 not
X70 VDD VSS DC_3 DC3 not
X71 VDD VSS DC_4 DC4 not
X72 VDD VSS DC_5 DC5 not
X73 VDD VSS DC_6 DC6 not
X74 VDD VSS DC_7 DC7 not
X75 VDD VSS DC_8 DC8 not
X76 VDD VSS DC_9 DC9 not
X77 VDD VSS DC_10 DC10 not
X78 VDD VSS DC_11 DC11 not
X79 VDD VSS DC_12 DC12 not
X80 VDD VSS DC_13 DC13 not
X81 VDD VSS DC_14 DC14 not
X82 VDD VSS DC_15 DC15 not
X83 VDD VSS DC_16 DC16 not
X84 VDD VSS DC_17 DC17 not
X85 VDD VSS DC_18 DC18 not
X86 VDD VSS DC_19 DC19 not
X87 VDD VSS DC_20 DC20 not
X88 VDD VSS DC_21 DC21 not
X89 VDD VSS DC_22 DC22 not
X90 VDD VSS DC_23 DC23 not
X91 VDD VSS DC_24 DC24 not
X92 VDD VSS DC_25 DC25 not
X93 VDD VSS DC_26 DC26 not
X94 VDD VSS DC_27 DC27 not
X95 VDD VSS DC_28 DC28 not
X96 VDD VSS DC_29 DC29 not
X97 VDD VSS DC_30 DC30 not
X98 VDD VSS DC_31 DC31 not
X99 VDD VSS DC_32 DC32 not
X100 VDD VSS DC_33 DC33 not
X101 VDD VSS DC_34 DC34 not
X102 VDD VSS DC_35 DC35 not
X103 VDD VSS DC_36 DC36 not
X104 VDD VSS DC_37 DC37 not
X105 VDD VSS DC_38 DC38 not
X106 VDD VSS DC_39 DC39 not
X107 VDD VSS DC_40 DC40 not
X108 VDD VSS DC_41 DC41 not
X109 VDD VSS DC_42 DC42 not
X110 VDD VSS DC_43 DC43 not
X111 VDD VSS DC_44 DC44 not
X112 VDD VSS DC_45 DC45 not
X113 VDD VSS DC_46 DC46 not
X114 VDD VSS DC_47 DC47 not
X115 VDD VSS DC_48 DC48 not
X116 VDD VSS DC_49 DC49 not
X117 VDD VSS DC_50 DC50 not
X118 VDD VSS DC_51 DC51 not
X119 VDD VSS DC_52 DC52 not
X120 VDD VSS DC_53 DC53 not
X121 VDD VSS DC_54 DC54 not
X122 VDD VSS DC_55 DC55 not
X123 VDD VSS DC_56 DC56 not
X124 VDD VSS DC_57 DC57 not
X125 VDD VSS DC_58 DC58 not
X126 VDD VSS DC_59 DC59 not
X127 VDD VSS DC_60 DC60 not
X128 VDD VSS DC_61 DC61 not
X129 VDD VSS DC_62 DC62 not
X130 VDD VSS DC_63 DC63 not
.ends row_dec64

.subckt row_driver VDD VSS WLEN A B
X0 VDD VSS A WLEN net1 nand2
X1 B net1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X2 B net1 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
.ends row_driver

.subckt rd_arr_64 VDD VSS WLEN DC0 DC1 DC2 DC3 DC4 DC5 DC6 DC7 DC8 DC9 DC10 DC11 DC12 DC13 DC14 DC15 DC16 DC17 DC18 DC19 DC20 DC21 DC22 DC23 DC24 DC25 DC26 DC27 DC28 DC29 DC30 DC31 DC32 DC33 DC34 DC35 DC36 DC37 DC38 DC39 DC40 DC41 DC42 DC43 DC44 DC45 DC46 DC47 DC48 DC49 DC50 DC51 DC52 DC53 DC54 DC55 DC56 DC57 DC58 DC59 DC60 DC61 DC62 DC63 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 WL32 WL33 WL34 WL35 WL36 WL37 WL38 WL39 WL40 WL41 WL42 WL43 WL44 WL45 WL46 WL47 WL48 WL49 WL50 WL51 WL52 WL53 WL54 WL55 WL56 WL57 WL58 WL59 WL60 WL61 WL62 WL63
X0 VDD VSS WLEN DC0 WL0 row_driver
X1 VDD VSS WLEN DC1 WL1 row_driver
X2 VDD VSS WLEN DC2 WL2 row_driver
X3 VDD VSS WLEN DC3 WL3 row_driver
X4 VDD VSS WLEN DC4 WL4 row_driver
X5 VDD VSS WLEN DC5 WL5 row_driver
X6 VDD VSS WLEN DC6 WL6 row_driver
X7 VDD VSS WLEN DC7 WL7 row_driver
X8 VDD VSS WLEN DC8 WL8 row_driver
X9 VDD VSS WLEN DC9 WL9 row_driver
X10 VDD VSS WLEN DC10 WL10 row_driver
X11 VDD VSS WLEN DC11 WL11 row_driver
X12 VDD VSS WLEN DC12 WL12 row_driver
X13 VDD VSS WLEN DC13 WL13 row_driver
X14 VDD VSS WLEN DC14 WL14 row_driver
X15 VDD VSS WLEN DC15 WL15 row_driver
X16 VDD VSS WLEN DC16 WL16 row_driver
X17 VDD VSS WLEN DC17 WL17 row_driver
X18 VDD VSS WLEN DC18 WL18 row_driver
X19 VDD VSS WLEN DC19 WL19 row_driver
X20 VDD VSS WLEN DC20 WL20 row_driver
X21 VDD VSS WLEN DC21 WL21 row_driver
X22 VDD VSS WLEN DC22 WL22 row_driver
X23 VDD VSS WLEN DC23 WL23 row_driver
X24 VDD VSS WLEN DC24 WL24 row_driver
X25 VDD VSS WLEN DC25 WL25 row_driver
X26 VDD VSS WLEN DC26 WL26 row_driver
X27 VDD VSS WLEN DC27 WL27 row_driver
X28 VDD VSS WLEN DC28 WL28 row_driver
X29 VDD VSS WLEN DC29 WL29 row_driver
X30 VDD VSS WLEN DC30 WL30 row_driver
X31 VDD VSS WLEN DC31 WL31 row_driver
X32 VDD VSS WLEN DC32 WL32 row_driver
X33 VDD VSS WLEN DC33 WL33 row_driver
X34 VDD VSS WLEN DC34 WL34 row_driver
X35 VDD VSS WLEN DC35 WL35 row_driver
X36 VDD VSS WLEN DC36 WL36 row_driver
X37 VDD VSS WLEN DC37 WL37 row_driver
X38 VDD VSS WLEN DC38 WL38 row_driver
X39 VDD VSS WLEN DC39 WL39 row_driver
X40 VDD VSS WLEN DC40 WL40 row_driver
X41 VDD VSS WLEN DC41 WL41 row_driver
X42 VDD VSS WLEN DC42 WL42 row_driver
X43 VDD VSS WLEN DC43 WL43 row_driver
X44 VDD VSS WLEN DC44 WL44 row_driver
X45 VDD VSS WLEN DC45 WL45 row_driver
X46 VDD VSS WLEN DC46 WL46 row_driver
X47 VDD VSS WLEN DC47 WL47 row_driver
X48 VDD VSS WLEN DC48 WL48 row_driver
X49 VDD VSS WLEN DC49 WL49 row_driver
X50 VDD VSS WLEN DC50 WL50 row_driver
X51 VDD VSS WLEN DC51 WL51 row_driver
X52 VDD VSS WLEN DC52 WL52 row_driver
X53 VDD VSS WLEN DC53 WL53 row_driver
X54 VDD VSS WLEN DC54 WL54 row_driver
X55 VDD VSS WLEN DC55 WL55 row_driver
X56 VDD VSS WLEN DC56 WL56 row_driver
X57 VDD VSS WLEN DC57 WL57 row_driver
X58 VDD VSS WLEN DC58 WL58 row_driver
X59 VDD VSS WLEN DC59 WL59 row_driver
X60 VDD VSS WLEN DC60 WL60 row_driver
X61 VDD VSS WLEN DC61 WL61 row_driver
X62 VDD VSS WLEN DC62 WL62 row_driver
X63 VDD VSS WLEN DC63 WL63 row_driver
.ends rd_arr_64

.subckt rd_arr_4 VDD VSS WLEN DC0 DC1 DC2 DC3 WL0 WL1 WL2 WL3
X0 VDD VSS WLEN DC0 WL0 row_driver
X1 VDD VSS WLEN DC1 WL1 row_driver
X2 VDD VSS WLEN DC2 WL2 row_driver
X3 VDD VSS WLEN DC3 WL3 row_driver
.ends rd_arr_4

.subckt col_dec4 VDD VSS A0 A1 DC0 DC1 DC2 DC3
X0 VDD VSS A1 A0 Y0 Y1 Y2 Y3 dec_2to4
X1 VDD VSS Y0 DC0 not
X2 VDD VSS Y1 DC1 not
X3 VDD VSS Y2 DC2 not
X4 VDD VSS Y3 DC3 not
.ends col_dec4

.subckt dido VDD VSS PCHG WREN SEL BL BL_ DW DW_ DR DR_
X0 BL_ net6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 BL net6 BL_ VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 BL net6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 net6 net5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 net6 net5 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X5 net5 PCHG VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X6 net5 PCHG VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X7 BL_ net4 DR_ VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X8 DR net4 BL VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X9 net4 SEL VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X10 BL net2 DW VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X11 DW_ net2 BL_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X12 net4 SEL VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X13 net3 net4 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X14 net3 net4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X15 VDD VSS net3 WREN net1 nand2
X16 VDD VSS net1 net2 not
.ends dido

.subckt dido_arr_128 VDD VSS PCHG WREN SEL0 SEL1 SEL2 SEL3 SEL4 SEL5 SEL6 SEL7 SEL8 SEL9 SEL10 SEL11 SEL12 SEL13 SEL14 SEL15 SEL16 SEL17 SEL18 SEL19 SEL20 SEL21 SEL22 SEL23 SEL24 SEL25 SEL26 SEL27 SEL28 SEL29 SEL30 SEL31 SEL32 SEL33 SEL34 SEL35 SEL36 SEL37 SEL38 SEL39 SEL40 SEL41 SEL42 SEL43 SEL44 SEL45 SEL46 SEL47 SEL48 SEL49 SEL50 SEL51 SEL52 SEL53 SEL54 SEL55 SEL56 SEL57 SEL58 SEL59 SEL60 SEL61 SEL62 SEL63 SEL64 SEL65 SEL66 SEL67 SEL68 SEL69 SEL70 SEL71 SEL72 SEL73 SEL74 SEL75 SEL76 SEL77 SEL78 SEL79 SEL80 SEL81 SEL82 SEL83 SEL84 SEL85 SEL86 SEL87 SEL88 SEL89 SEL90 SEL91 SEL92 SEL93 SEL94 SEL95 SEL96 SEL97 SEL98 SEL99 SEL100 SEL101 SEL102 SEL103 SEL104 SEL105 SEL106 SEL107 SEL108 SEL109 SEL110 SEL111 SEL112 SEL113 SEL114 SEL115 SEL116 SEL117 SEL118 SEL119 SEL120 SEL121 SEL122 SEL123 SEL124 SEL125 SEL126 SEL127 BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 DW0 DW_0 DW1 DW_1 DW2 DW_2 DW3 DW_3 DW4 DW_4 DW5 DW_5 DW6 DW_6 DW7 DW_7 DW8 DW_8 DW9 DW_9 DW10 DW_10 DW11 DW_11 DW12 DW_12 DW13 DW_13 DW14 DW_14 DW15 DW_15 DW16 DW_16 DW17 DW_17 DW18 DW_18 DW19 DW_19 DW20 DW_20 DW21 DW_21 DW22 DW_22 DW23 DW_23 DW24 DW_24 DW25 DW_25 DW26 DW_26 DW27 DW_27 DW28 DW_28 DW29 DW_29 DW30 DW_30 DW31 DW_31 DW32 DW_32 DW33 DW_33 DW34 DW_34 DW35 DW_35 DW36 DW_36 DW37 DW_37 DW38 DW_38 DW39 DW_39 DW40 DW_40 DW41 DW_41 DW42 DW_42 DW43 DW_43 DW44 DW_44 DW45 DW_45 DW46 DW_46 DW47 DW_47 DW48 DW_48 DW49 DW_49 DW50 DW_50 DW51 DW_51 DW52 DW_52 DW53 DW_53 DW54 DW_54 DW55 DW_55 DW56 DW_56 DW57 DW_57 DW58 DW_58 DW59 DW_59 DW60 DW_60 DW61 DW_61 DW62 DW_62 DW63 DW_63 DW64 DW_64 DW65 DW_65 DW66 DW_66 DW67 DW_67 DW68 DW_68 DW69 DW_69 DW70 DW_70 DW71 DW_71 DW72 DW_72 DW73 DW_73 DW74 DW_74 DW75 DW_75 DW76 DW_76 DW77 DW_77 DW78 DW_78 DW79 DW_79 DW80 DW_80 DW81 DW_81 DW82 DW_82 DW83 DW_83 DW84 DW_84 DW85 DW_85 DW86 DW_86 DW87 DW_87 DW88 DW_88 DW89 DW_89 DW90 DW_90 DW91 DW_91 DW92 DW_92 DW93 DW_93 DW94 DW_94 DW95 DW_95 DW96 DW_96 DW97 DW_97 DW98 DW_98 DW99 DW_99 DW100 DW_100 DW101 DW_101 DW102 DW_102 DW103 DW_103 DW104 DW_104 DW105 DW_105 DW106 DW_106 DW107 DW_107 DW108 DW_108 DW109 DW_109 DW110 DW_110 DW111 DW_111 DW112 DW_112 DW113 DW_113 DW114 DW_114 DW115 DW_115 DW116 DW_116 DW117 DW_117 DW118 DW_118 DW119 DW_119 DW120 DW_120 DW121 DW_121 DW122 DW_122 DW123 DW_123 DW124 DW_124 DW125 DW_125 DW126 DW_126 DW127 DW_127 DR0 DR_0 DR1 DR_1 DR2 DR_2 DR3 DR_3 DR4 DR_4 DR5 DR_5 DR6 DR_6 DR7 DR_7 DR8 DR_8 DR9 DR_9 DR10 DR_10 DR11 DR_11 DR12 DR_12 DR13 DR_13 DR14 DR_14 DR15 DR_15 DR16 DR_16 DR17 DR_17 DR18 DR_18 DR19 DR_19 DR20 DR_20 DR21 DR_21 DR22 DR_22 DR23 DR_23 DR24 DR_24 DR25 DR_25 DR26 DR_26 DR27 DR_27 DR28 DR_28 DR29 DR_29 DR30 DR_30 DR31 DR_31 DR32 DR_32 DR33 DR_33 DR34 DR_34 DR35 DR_35 DR36 DR_36 DR37 DR_37 DR38 DR_38 DR39 DR_39 DR40 DR_40 DR41 DR_41 DR42 DR_42 DR43 DR_43 DR44 DR_44 DR45 DR_45 DR46 DR_46 DR47 DR_47 DR48 DR_48 DR49 DR_49 DR50 DR_50 DR51 DR_51 DR52 DR_52 DR53 DR_53 DR54 DR_54 DR55 DR_55 DR56 DR_56 DR57 DR_57 DR58 DR_58 DR59 DR_59 DR60 DR_60 DR61 DR_61 DR62 DR_62 DR63 DR_63 DR64 DR_64 DR65 DR_65 DR66 DR_66 DR67 DR_67 DR68 DR_68 DR69 DR_69 DR70 DR_70 DR71 DR_71 DR72 DR_72 DR73 DR_73 DR74 DR_74 DR75 DR_75 DR76 DR_76 DR77 DR_77 DR78 DR_78 DR79 DR_79 DR80 DR_80 DR81 DR_81 DR82 DR_82 DR83 DR_83 DR84 DR_84 DR85 DR_85 DR86 DR_86 DR87 DR_87 DR88 DR_88 DR89 DR_89 DR90 DR_90 DR91 DR_91 DR92 DR_92 DR93 DR_93 DR94 DR_94 DR95 DR_95 DR96 DR_96 DR97 DR_97 DR98 DR_98 DR99 DR_99 DR100 DR_100 DR101 DR_101 DR102 DR_102 DR103 DR_103 DR104 DR_104 DR105 DR_105 DR106 DR_106 DR107 DR_107 DR108 DR_108 DR109 DR_109 DR110 DR_110 DR111 DR_111 DR112 DR_112 DR113 DR_113 DR114 DR_114 DR115 DR_115 DR116 DR_116 DR117 DR_117 DR118 DR_118 DR119 DR_119 DR120 DR_120 DR121 DR_121 DR122 DR_122 DR123 DR_123 DR124 DR_124 DR125 DR_125 DR126 DR_126 DR127 DR_127
X0 VDD VSS PCHG WREN SEL0 BL0 BL_0 DW0 DW_0 DR0 DR_0 dido
X1 VDD VSS PCHG WREN SEL1 BL1 BL_1 DW1 DW_1 DR1 DR_1 dido
X2 VDD VSS PCHG WREN SEL2 BL2 BL_2 DW2 DW_2 DR2 DR_2 dido
X3 VDD VSS PCHG WREN SEL3 BL3 BL_3 DW3 DW_3 DR3 DR_3 dido
X4 VDD VSS PCHG WREN SEL4 BL4 BL_4 DW4 DW_4 DR4 DR_4 dido
X5 VDD VSS PCHG WREN SEL5 BL5 BL_5 DW5 DW_5 DR5 DR_5 dido
X6 VDD VSS PCHG WREN SEL6 BL6 BL_6 DW6 DW_6 DR6 DR_6 dido
X7 VDD VSS PCHG WREN SEL7 BL7 BL_7 DW7 DW_7 DR7 DR_7 dido
X8 VDD VSS PCHG WREN SEL8 BL8 BL_8 DW8 DW_8 DR8 DR_8 dido
X9 VDD VSS PCHG WREN SEL9 BL9 BL_9 DW9 DW_9 DR9 DR_9 dido
X10 VDD VSS PCHG WREN SEL10 BL10 BL_10 DW10 DW_10 DR10 DR_10 dido
X11 VDD VSS PCHG WREN SEL11 BL11 BL_11 DW11 DW_11 DR11 DR_11 dido
X12 VDD VSS PCHG WREN SEL12 BL12 BL_12 DW12 DW_12 DR12 DR_12 dido
X13 VDD VSS PCHG WREN SEL13 BL13 BL_13 DW13 DW_13 DR13 DR_13 dido
X14 VDD VSS PCHG WREN SEL14 BL14 BL_14 DW14 DW_14 DR14 DR_14 dido
X15 VDD VSS PCHG WREN SEL15 BL15 BL_15 DW15 DW_15 DR15 DR_15 dido
X16 VDD VSS PCHG WREN SEL16 BL16 BL_16 DW16 DW_16 DR16 DR_16 dido
X17 VDD VSS PCHG WREN SEL17 BL17 BL_17 DW17 DW_17 DR17 DR_17 dido
X18 VDD VSS PCHG WREN SEL18 BL18 BL_18 DW18 DW_18 DR18 DR_18 dido
X19 VDD VSS PCHG WREN SEL19 BL19 BL_19 DW19 DW_19 DR19 DR_19 dido
X20 VDD VSS PCHG WREN SEL20 BL20 BL_20 DW20 DW_20 DR20 DR_20 dido
X21 VDD VSS PCHG WREN SEL21 BL21 BL_21 DW21 DW_21 DR21 DR_21 dido
X22 VDD VSS PCHG WREN SEL22 BL22 BL_22 DW22 DW_22 DR22 DR_22 dido
X23 VDD VSS PCHG WREN SEL23 BL23 BL_23 DW23 DW_23 DR23 DR_23 dido
X24 VDD VSS PCHG WREN SEL24 BL24 BL_24 DW24 DW_24 DR24 DR_24 dido
X25 VDD VSS PCHG WREN SEL25 BL25 BL_25 DW25 DW_25 DR25 DR_25 dido
X26 VDD VSS PCHG WREN SEL26 BL26 BL_26 DW26 DW_26 DR26 DR_26 dido
X27 VDD VSS PCHG WREN SEL27 BL27 BL_27 DW27 DW_27 DR27 DR_27 dido
X28 VDD VSS PCHG WREN SEL28 BL28 BL_28 DW28 DW_28 DR28 DR_28 dido
X29 VDD VSS PCHG WREN SEL29 BL29 BL_29 DW29 DW_29 DR29 DR_29 dido
X30 VDD VSS PCHG WREN SEL30 BL30 BL_30 DW30 DW_30 DR30 DR_30 dido
X31 VDD VSS PCHG WREN SEL31 BL31 BL_31 DW31 DW_31 DR31 DR_31 dido
X32 VDD VSS PCHG WREN SEL32 BL32 BL_32 DW32 DW_32 DR32 DR_32 dido
X33 VDD VSS PCHG WREN SEL33 BL33 BL_33 DW33 DW_33 DR33 DR_33 dido
X34 VDD VSS PCHG WREN SEL34 BL34 BL_34 DW34 DW_34 DR34 DR_34 dido
X35 VDD VSS PCHG WREN SEL35 BL35 BL_35 DW35 DW_35 DR35 DR_35 dido
X36 VDD VSS PCHG WREN SEL36 BL36 BL_36 DW36 DW_36 DR36 DR_36 dido
X37 VDD VSS PCHG WREN SEL37 BL37 BL_37 DW37 DW_37 DR37 DR_37 dido
X38 VDD VSS PCHG WREN SEL38 BL38 BL_38 DW38 DW_38 DR38 DR_38 dido
X39 VDD VSS PCHG WREN SEL39 BL39 BL_39 DW39 DW_39 DR39 DR_39 dido
X40 VDD VSS PCHG WREN SEL40 BL40 BL_40 DW40 DW_40 DR40 DR_40 dido
X41 VDD VSS PCHG WREN SEL41 BL41 BL_41 DW41 DW_41 DR41 DR_41 dido
X42 VDD VSS PCHG WREN SEL42 BL42 BL_42 DW42 DW_42 DR42 DR_42 dido
X43 VDD VSS PCHG WREN SEL43 BL43 BL_43 DW43 DW_43 DR43 DR_43 dido
X44 VDD VSS PCHG WREN SEL44 BL44 BL_44 DW44 DW_44 DR44 DR_44 dido
X45 VDD VSS PCHG WREN SEL45 BL45 BL_45 DW45 DW_45 DR45 DR_45 dido
X46 VDD VSS PCHG WREN SEL46 BL46 BL_46 DW46 DW_46 DR46 DR_46 dido
X47 VDD VSS PCHG WREN SEL47 BL47 BL_47 DW47 DW_47 DR47 DR_47 dido
X48 VDD VSS PCHG WREN SEL48 BL48 BL_48 DW48 DW_48 DR48 DR_48 dido
X49 VDD VSS PCHG WREN SEL49 BL49 BL_49 DW49 DW_49 DR49 DR_49 dido
X50 VDD VSS PCHG WREN SEL50 BL50 BL_50 DW50 DW_50 DR50 DR_50 dido
X51 VDD VSS PCHG WREN SEL51 BL51 BL_51 DW51 DW_51 DR51 DR_51 dido
X52 VDD VSS PCHG WREN SEL52 BL52 BL_52 DW52 DW_52 DR52 DR_52 dido
X53 VDD VSS PCHG WREN SEL53 BL53 BL_53 DW53 DW_53 DR53 DR_53 dido
X54 VDD VSS PCHG WREN SEL54 BL54 BL_54 DW54 DW_54 DR54 DR_54 dido
X55 VDD VSS PCHG WREN SEL55 BL55 BL_55 DW55 DW_55 DR55 DR_55 dido
X56 VDD VSS PCHG WREN SEL56 BL56 BL_56 DW56 DW_56 DR56 DR_56 dido
X57 VDD VSS PCHG WREN SEL57 BL57 BL_57 DW57 DW_57 DR57 DR_57 dido
X58 VDD VSS PCHG WREN SEL58 BL58 BL_58 DW58 DW_58 DR58 DR_58 dido
X59 VDD VSS PCHG WREN SEL59 BL59 BL_59 DW59 DW_59 DR59 DR_59 dido
X60 VDD VSS PCHG WREN SEL60 BL60 BL_60 DW60 DW_60 DR60 DR_60 dido
X61 VDD VSS PCHG WREN SEL61 BL61 BL_61 DW61 DW_61 DR61 DR_61 dido
X62 VDD VSS PCHG WREN SEL62 BL62 BL_62 DW62 DW_62 DR62 DR_62 dido
X63 VDD VSS PCHG WREN SEL63 BL63 BL_63 DW63 DW_63 DR63 DR_63 dido
X64 VDD VSS PCHG WREN SEL64 BL64 BL_64 DW64 DW_64 DR64 DR_64 dido
X65 VDD VSS PCHG WREN SEL65 BL65 BL_65 DW65 DW_65 DR65 DR_65 dido
X66 VDD VSS PCHG WREN SEL66 BL66 BL_66 DW66 DW_66 DR66 DR_66 dido
X67 VDD VSS PCHG WREN SEL67 BL67 BL_67 DW67 DW_67 DR67 DR_67 dido
X68 VDD VSS PCHG WREN SEL68 BL68 BL_68 DW68 DW_68 DR68 DR_68 dido
X69 VDD VSS PCHG WREN SEL69 BL69 BL_69 DW69 DW_69 DR69 DR_69 dido
X70 VDD VSS PCHG WREN SEL70 BL70 BL_70 DW70 DW_70 DR70 DR_70 dido
X71 VDD VSS PCHG WREN SEL71 BL71 BL_71 DW71 DW_71 DR71 DR_71 dido
X72 VDD VSS PCHG WREN SEL72 BL72 BL_72 DW72 DW_72 DR72 DR_72 dido
X73 VDD VSS PCHG WREN SEL73 BL73 BL_73 DW73 DW_73 DR73 DR_73 dido
X74 VDD VSS PCHG WREN SEL74 BL74 BL_74 DW74 DW_74 DR74 DR_74 dido
X75 VDD VSS PCHG WREN SEL75 BL75 BL_75 DW75 DW_75 DR75 DR_75 dido
X76 VDD VSS PCHG WREN SEL76 BL76 BL_76 DW76 DW_76 DR76 DR_76 dido
X77 VDD VSS PCHG WREN SEL77 BL77 BL_77 DW77 DW_77 DR77 DR_77 dido
X78 VDD VSS PCHG WREN SEL78 BL78 BL_78 DW78 DW_78 DR78 DR_78 dido
X79 VDD VSS PCHG WREN SEL79 BL79 BL_79 DW79 DW_79 DR79 DR_79 dido
X80 VDD VSS PCHG WREN SEL80 BL80 BL_80 DW80 DW_80 DR80 DR_80 dido
X81 VDD VSS PCHG WREN SEL81 BL81 BL_81 DW81 DW_81 DR81 DR_81 dido
X82 VDD VSS PCHG WREN SEL82 BL82 BL_82 DW82 DW_82 DR82 DR_82 dido
X83 VDD VSS PCHG WREN SEL83 BL83 BL_83 DW83 DW_83 DR83 DR_83 dido
X84 VDD VSS PCHG WREN SEL84 BL84 BL_84 DW84 DW_84 DR84 DR_84 dido
X85 VDD VSS PCHG WREN SEL85 BL85 BL_85 DW85 DW_85 DR85 DR_85 dido
X86 VDD VSS PCHG WREN SEL86 BL86 BL_86 DW86 DW_86 DR86 DR_86 dido
X87 VDD VSS PCHG WREN SEL87 BL87 BL_87 DW87 DW_87 DR87 DR_87 dido
X88 VDD VSS PCHG WREN SEL88 BL88 BL_88 DW88 DW_88 DR88 DR_88 dido
X89 VDD VSS PCHG WREN SEL89 BL89 BL_89 DW89 DW_89 DR89 DR_89 dido
X90 VDD VSS PCHG WREN SEL90 BL90 BL_90 DW90 DW_90 DR90 DR_90 dido
X91 VDD VSS PCHG WREN SEL91 BL91 BL_91 DW91 DW_91 DR91 DR_91 dido
X92 VDD VSS PCHG WREN SEL92 BL92 BL_92 DW92 DW_92 DR92 DR_92 dido
X93 VDD VSS PCHG WREN SEL93 BL93 BL_93 DW93 DW_93 DR93 DR_93 dido
X94 VDD VSS PCHG WREN SEL94 BL94 BL_94 DW94 DW_94 DR94 DR_94 dido
X95 VDD VSS PCHG WREN SEL95 BL95 BL_95 DW95 DW_95 DR95 DR_95 dido
X96 VDD VSS PCHG WREN SEL96 BL96 BL_96 DW96 DW_96 DR96 DR_96 dido
X97 VDD VSS PCHG WREN SEL97 BL97 BL_97 DW97 DW_97 DR97 DR_97 dido
X98 VDD VSS PCHG WREN SEL98 BL98 BL_98 DW98 DW_98 DR98 DR_98 dido
X99 VDD VSS PCHG WREN SEL99 BL99 BL_99 DW99 DW_99 DR99 DR_99 dido
X100 VDD VSS PCHG WREN SEL100 BL100 BL_100 DW100 DW_100 DR100 DR_100 dido
X101 VDD VSS PCHG WREN SEL101 BL101 BL_101 DW101 DW_101 DR101 DR_101 dido
X102 VDD VSS PCHG WREN SEL102 BL102 BL_102 DW102 DW_102 DR102 DR_102 dido
X103 VDD VSS PCHG WREN SEL103 BL103 BL_103 DW103 DW_103 DR103 DR_103 dido
X104 VDD VSS PCHG WREN SEL104 BL104 BL_104 DW104 DW_104 DR104 DR_104 dido
X105 VDD VSS PCHG WREN SEL105 BL105 BL_105 DW105 DW_105 DR105 DR_105 dido
X106 VDD VSS PCHG WREN SEL106 BL106 BL_106 DW106 DW_106 DR106 DR_106 dido
X107 VDD VSS PCHG WREN SEL107 BL107 BL_107 DW107 DW_107 DR107 DR_107 dido
X108 VDD VSS PCHG WREN SEL108 BL108 BL_108 DW108 DW_108 DR108 DR_108 dido
X109 VDD VSS PCHG WREN SEL109 BL109 BL_109 DW109 DW_109 DR109 DR_109 dido
X110 VDD VSS PCHG WREN SEL110 BL110 BL_110 DW110 DW_110 DR110 DR_110 dido
X111 VDD VSS PCHG WREN SEL111 BL111 BL_111 DW111 DW_111 DR111 DR_111 dido
X112 VDD VSS PCHG WREN SEL112 BL112 BL_112 DW112 DW_112 DR112 DR_112 dido
X113 VDD VSS PCHG WREN SEL113 BL113 BL_113 DW113 DW_113 DR113 DR_113 dido
X114 VDD VSS PCHG WREN SEL114 BL114 BL_114 DW114 DW_114 DR114 DR_114 dido
X115 VDD VSS PCHG WREN SEL115 BL115 BL_115 DW115 DW_115 DR115 DR_115 dido
X116 VDD VSS PCHG WREN SEL116 BL116 BL_116 DW116 DW_116 DR116 DR_116 dido
X117 VDD VSS PCHG WREN SEL117 BL117 BL_117 DW117 DW_117 DR117 DR_117 dido
X118 VDD VSS PCHG WREN SEL118 BL118 BL_118 DW118 DW_118 DR118 DR_118 dido
X119 VDD VSS PCHG WREN SEL119 BL119 BL_119 DW119 DW_119 DR119 DR_119 dido
X120 VDD VSS PCHG WREN SEL120 BL120 BL_120 DW120 DW_120 DR120 DR_120 dido
X121 VDD VSS PCHG WREN SEL121 BL121 BL_121 DW121 DW_121 DR121 DR_121 dido
X122 VDD VSS PCHG WREN SEL122 BL122 BL_122 DW122 DW_122 DR122 DR_122 dido
X123 VDD VSS PCHG WREN SEL123 BL123 BL_123 DW123 DW_123 DR123 DR_123 dido
X124 VDD VSS PCHG WREN SEL124 BL124 BL_124 DW124 DW_124 DR124 DR_124 dido
X125 VDD VSS PCHG WREN SEL125 BL125 BL_125 DW125 DW_125 DR125 DR_125 dido
X126 VDD VSS PCHG WREN SEL126 BL126 BL_126 DW126 DW_126 DR126 DR_126 dido
X127 VDD VSS PCHG WREN SEL127 BL127 BL_127 DW127 DW_127 DR127 DR_127 dido
.ends dido_arr_128

.subckt write_driver VDD VSS WREN Din DW DW_
X0 en_ WREN VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 en_ WREN VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X4 d_ Din VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X5 d_ Din VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X6 net1 Din VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X7 DW_ en_ net1 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X8 DW_ WREN net2 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
X9 net2 Din VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
X10 net3 d_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X11 DW en_ net3 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X12 DW WREN net4 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
X13 net4 d_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
.ends write_driver

.subckt del10 VDD VSS A B
X0 VDD VSS A net1 notdel
X1 VDD VSS net1 net2 notdel
X2 VDD VSS net2 net3 notdel
X3 VDD VSS net3 net4 notdel
X4 VDD VSS net4 net5 notdel
X5 VDD VSS net5 net6 notdel
X6 VDD VSS net6 net7 notdel
X7 VDD VSS net7 net8 notdel
X8 VDD VSS net8 net9 notdel
X9 VDD VSS net9 net10 notdel
X10 VDD VSS net10 net11 notdel
X11 VDD VSS A net11 net12 nand2
X12 VDD VSS net12 B not
.ends del10

.subckt ctrl VDD VSS clk cs write DBL DBL_ WREN PCHG WLEN SAEN
X0 clk_ clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 clk_ clk VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X2 WLENP clk_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 WLENP clk_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X4 VDD VSS write WREN_ not
X8 PCHG clk_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X9 PCHG clk_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
X10 DBL_ PCHG VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X11 DBL PCHG DBL_ VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X12 DBL PCHG VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X13 VDD VSS cs WLENP WLENPP nand2
X21 WLEN WLENPP VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X22 WLEN WLENPP VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
X15 VDD VSS DBL_ RBL not
X16 VDD VSS WLEN RBL SAEN_ nand2
X17 SAEN SAEN_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X18 SAEN SAEN_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
X19 WREN WREN_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X20 WREN WREN_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
.ends ctrl

.subckt input_reg9 VDD VSS clk D0 D1 D2 D3 D4 D5 D6 D7 D8 Q0 Q1 Q2 Q3 Q4 Q5 Q6 Q7 Q8
X0 VDD VSS clk D0 Q0 in_reg
X1 VDD VSS clk D1 Q1 in_reg
X2 VDD VSS clk D2 Q2 in_reg
X3 VDD VSS clk D3 Q3 in_reg
X4 VDD VSS clk D4 Q4 in_reg
X5 VDD VSS clk D5 Q5 in_reg
X6 VDD VSS clk D6 Q6 in_reg
X7 VDD VSS clk D7 Q7 in_reg
X8 VDD VSS clk D8 Q8 in_reg
.ends input_reg9

.subckt datain_reg32 VDD VSS clk WREN din0 din1 din2 din3 din4 din5 din6 din7 din8 din9 din10 din11 din12 din13 din14 din15 din16 din17 din18 din19 din20 din21 din22 din23 din24 din25 din26 din27 din28 din29 din30 din31 DW0 DW_0 DW1 DW_1 DW2 DW_2 DW3 DW_3 DW4 DW_4 DW5 DW_5 DW6 DW_6 DW7 DW_7 DW8 DW_8 DW9 DW_9 DW10 DW_10 DW11 DW_11 DW12 DW_12 DW13 DW_13 DW14 DW_14 DW15 DW_15 DW16 DW_16 DW17 DW_17 DW18 DW_18 DW19 DW_19 DW20 DW_20 DW21 DW_21 DW22 DW_22 DW23 DW_23 DW24 DW_24 DW25 DW_25 DW26 DW_26 DW27 DW_27 DW28 DW_28 DW29 DW_29 DW30 DW_30 DW31 DW_31
X0 VDD VSS clk din0 din_r0 in_reg
X1 VDD VSS clk din1 din_r1 in_reg
X2 VDD VSS clk din2 din_r2 in_reg
X3 VDD VSS clk din3 din_r3 in_reg
X4 VDD VSS clk din4 din_r4 in_reg
X5 VDD VSS clk din5 din_r5 in_reg
X6 VDD VSS clk din6 din_r6 in_reg
X7 VDD VSS clk din7 din_r7 in_reg
X8 VDD VSS clk din8 din_r8 in_reg
X9 VDD VSS clk din9 din_r9 in_reg
X10 VDD VSS clk din10 din_r10 in_reg
X11 VDD VSS clk din11 din_r11 in_reg
X12 VDD VSS clk din12 din_r12 in_reg
X13 VDD VSS clk din13 din_r13 in_reg
X14 VDD VSS clk din14 din_r14 in_reg
X15 VDD VSS clk din15 din_r15 in_reg
X16 VDD VSS clk din16 din_r16 in_reg
X17 VDD VSS clk din17 din_r17 in_reg
X18 VDD VSS clk din18 din_r18 in_reg
X19 VDD VSS clk din19 din_r19 in_reg
X20 VDD VSS clk din20 din_r20 in_reg
X21 VDD VSS clk din21 din_r21 in_reg
X22 VDD VSS clk din22 din_r22 in_reg
X23 VDD VSS clk din23 din_r23 in_reg
X24 VDD VSS clk din24 din_r24 in_reg
X25 VDD VSS clk din25 din_r25 in_reg
X26 VDD VSS clk din26 din_r26 in_reg
X27 VDD VSS clk din27 din_r27 in_reg
X28 VDD VSS clk din28 din_r28 in_reg
X29 VDD VSS clk din29 din_r29 in_reg
X30 VDD VSS clk din30 din_r30 in_reg
X31 VDD VSS clk din31 din_r31 in_reg
X32 VDD VSS WREN din_r0 DW0 DW_0 write_driver
X36 VDD VSS WREN din_r1 DW1 DW_1 write_driver
X40 VDD VSS WREN din_r2 DW2 DW_2 write_driver
X44 VDD VSS WREN din_r3 DW3 DW_3 write_driver
X48 VDD VSS WREN din_r4 DW4 DW_4 write_driver
X52 VDD VSS WREN din_r5 DW5 DW_5 write_driver
X56 VDD VSS WREN din_r6 DW6 DW_6 write_driver
X60 VDD VSS WREN din_r7 DW7 DW_7 write_driver
X64 VDD VSS WREN din_r8 DW8 DW_8 write_driver
X68 VDD VSS WREN din_r9 DW9 DW_9 write_driver
X72 VDD VSS WREN din_r10 DW10 DW_10 write_driver
X76 VDD VSS WREN din_r11 DW11 DW_11 write_driver
X80 VDD VSS WREN din_r12 DW12 DW_12 write_driver
X84 VDD VSS WREN din_r13 DW13 DW_13 write_driver
X88 VDD VSS WREN din_r14 DW14 DW_14 write_driver
X92 VDD VSS WREN din_r15 DW15 DW_15 write_driver
X96 VDD VSS WREN din_r16 DW16 DW_16 write_driver
X100 VDD VSS WREN din_r17 DW17 DW_17 write_driver
X104 VDD VSS WREN din_r18 DW18 DW_18 write_driver
X108 VDD VSS WREN din_r19 DW19 DW_19 write_driver
X112 VDD VSS WREN din_r20 DW20 DW_20 write_driver
X116 VDD VSS WREN din_r21 DW21 DW_21 write_driver
X120 VDD VSS WREN din_r22 DW22 DW_22 write_driver
X124 VDD VSS WREN din_r23 DW23 DW_23 write_driver
X128 VDD VSS WREN din_r24 DW24 DW_24 write_driver
X132 VDD VSS WREN din_r25 DW25 DW_25 write_driver
X136 VDD VSS WREN din_r26 DW26 DW_26 write_driver
X140 VDD VSS WREN din_r27 DW27 DW_27 write_driver
X144 VDD VSS WREN din_r28 DW28 DW_28 write_driver
X148 VDD VSS WREN din_r29 DW29 DW_29 write_driver
X152 VDD VSS WREN din_r30 DW30 DW_30 write_driver
X156 VDD VSS WREN din_r31 DW31 DW_31 write_driver
.ends datain_reg32

.subckt bit_arr_128 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL
X0 VDD VSS WL BL0 BL_0 bit_cell
X1 VDD VSS WL BL1 BL_1 bit_cell
X2 VDD VSS WL BL2 BL_2 bit_cell
X3 VDD VSS WL BL3 BL_3 bit_cell
X4 VDD VSS WL BL4 BL_4 bit_cell
X5 VDD VSS WL BL5 BL_5 bit_cell
X6 VDD VSS WL BL6 BL_6 bit_cell
X7 VDD VSS WL BL7 BL_7 bit_cell
X8 VDD VSS WL BL8 BL_8 bit_cell
X9 VDD VSS WL BL9 BL_9 bit_cell
X10 VDD VSS WL BL10 BL_10 bit_cell
X11 VDD VSS WL BL11 BL_11 bit_cell
X12 VDD VSS WL BL12 BL_12 bit_cell
X13 VDD VSS WL BL13 BL_13 bit_cell
X14 VDD VSS WL BL14 BL_14 bit_cell
X15 VDD VSS WL BL15 BL_15 bit_cell
X16 VDD VSS WL BL16 BL_16 bit_cell
X17 VDD VSS WL BL17 BL_17 bit_cell
X18 VDD VSS WL BL18 BL_18 bit_cell
X19 VDD VSS WL BL19 BL_19 bit_cell
X20 VDD VSS WL BL20 BL_20 bit_cell
X21 VDD VSS WL BL21 BL_21 bit_cell
X22 VDD VSS WL BL22 BL_22 bit_cell
X23 VDD VSS WL BL23 BL_23 bit_cell
X24 VDD VSS WL BL24 BL_24 bit_cell
X25 VDD VSS WL BL25 BL_25 bit_cell
X26 VDD VSS WL BL26 BL_26 bit_cell
X27 VDD VSS WL BL27 BL_27 bit_cell
X28 VDD VSS WL BL28 BL_28 bit_cell
X29 VDD VSS WL BL29 BL_29 bit_cell
X30 VDD VSS WL BL30 BL_30 bit_cell
X31 VDD VSS WL BL31 BL_31 bit_cell
X32 VDD VSS WL BL32 BL_32 bit_cell
X33 VDD VSS WL BL33 BL_33 bit_cell
X34 VDD VSS WL BL34 BL_34 bit_cell
X35 VDD VSS WL BL35 BL_35 bit_cell
X36 VDD VSS WL BL36 BL_36 bit_cell
X37 VDD VSS WL BL37 BL_37 bit_cell
X38 VDD VSS WL BL38 BL_38 bit_cell
X39 VDD VSS WL BL39 BL_39 bit_cell
X40 VDD VSS WL BL40 BL_40 bit_cell
X41 VDD VSS WL BL41 BL_41 bit_cell
X42 VDD VSS WL BL42 BL_42 bit_cell
X43 VDD VSS WL BL43 BL_43 bit_cell
X44 VDD VSS WL BL44 BL_44 bit_cell
X45 VDD VSS WL BL45 BL_45 bit_cell
X46 VDD VSS WL BL46 BL_46 bit_cell
X47 VDD VSS WL BL47 BL_47 bit_cell
X48 VDD VSS WL BL48 BL_48 bit_cell
X49 VDD VSS WL BL49 BL_49 bit_cell
X50 VDD VSS WL BL50 BL_50 bit_cell
X51 VDD VSS WL BL51 BL_51 bit_cell
X52 VDD VSS WL BL52 BL_52 bit_cell
X53 VDD VSS WL BL53 BL_53 bit_cell
X54 VDD VSS WL BL54 BL_54 bit_cell
X55 VDD VSS WL BL55 BL_55 bit_cell
X56 VDD VSS WL BL56 BL_56 bit_cell
X57 VDD VSS WL BL57 BL_57 bit_cell
X58 VDD VSS WL BL58 BL_58 bit_cell
X59 VDD VSS WL BL59 BL_59 bit_cell
X60 VDD VSS WL BL60 BL_60 bit_cell
X61 VDD VSS WL BL61 BL_61 bit_cell
X62 VDD VSS WL BL62 BL_62 bit_cell
X63 VDD VSS WL BL63 BL_63 bit_cell
X64 VDD VSS WL BL64 BL_64 bit_cell
X65 VDD VSS WL BL65 BL_65 bit_cell
X66 VDD VSS WL BL66 BL_66 bit_cell
X67 VDD VSS WL BL67 BL_67 bit_cell
X68 VDD VSS WL BL68 BL_68 bit_cell
X69 VDD VSS WL BL69 BL_69 bit_cell
X70 VDD VSS WL BL70 BL_70 bit_cell
X71 VDD VSS WL BL71 BL_71 bit_cell
X72 VDD VSS WL BL72 BL_72 bit_cell
X73 VDD VSS WL BL73 BL_73 bit_cell
X74 VDD VSS WL BL74 BL_74 bit_cell
X75 VDD VSS WL BL75 BL_75 bit_cell
X76 VDD VSS WL BL76 BL_76 bit_cell
X77 VDD VSS WL BL77 BL_77 bit_cell
X78 VDD VSS WL BL78 BL_78 bit_cell
X79 VDD VSS WL BL79 BL_79 bit_cell
X80 VDD VSS WL BL80 BL_80 bit_cell
X81 VDD VSS WL BL81 BL_81 bit_cell
X82 VDD VSS WL BL82 BL_82 bit_cell
X83 VDD VSS WL BL83 BL_83 bit_cell
X84 VDD VSS WL BL84 BL_84 bit_cell
X85 VDD VSS WL BL85 BL_85 bit_cell
X86 VDD VSS WL BL86 BL_86 bit_cell
X87 VDD VSS WL BL87 BL_87 bit_cell
X88 VDD VSS WL BL88 BL_88 bit_cell
X89 VDD VSS WL BL89 BL_89 bit_cell
X90 VDD VSS WL BL90 BL_90 bit_cell
X91 VDD VSS WL BL91 BL_91 bit_cell
X92 VDD VSS WL BL92 BL_92 bit_cell
X93 VDD VSS WL BL93 BL_93 bit_cell
X94 VDD VSS WL BL94 BL_94 bit_cell
X95 VDD VSS WL BL95 BL_95 bit_cell
X96 VDD VSS WL BL96 BL_96 bit_cell
X97 VDD VSS WL BL97 BL_97 bit_cell
X98 VDD VSS WL BL98 BL_98 bit_cell
X99 VDD VSS WL BL99 BL_99 bit_cell
X100 VDD VSS WL BL100 BL_100 bit_cell
X101 VDD VSS WL BL101 BL_101 bit_cell
X102 VDD VSS WL BL102 BL_102 bit_cell
X103 VDD VSS WL BL103 BL_103 bit_cell
X104 VDD VSS WL BL104 BL_104 bit_cell
X105 VDD VSS WL BL105 BL_105 bit_cell
X106 VDD VSS WL BL106 BL_106 bit_cell
X107 VDD VSS WL BL107 BL_107 bit_cell
X108 VDD VSS WL BL108 BL_108 bit_cell
X109 VDD VSS WL BL109 BL_109 bit_cell
X110 VDD VSS WL BL110 BL_110 bit_cell
X111 VDD VSS WL BL111 BL_111 bit_cell
X112 VDD VSS WL BL112 BL_112 bit_cell
X113 VDD VSS WL BL113 BL_113 bit_cell
X114 VDD VSS WL BL114 BL_114 bit_cell
X115 VDD VSS WL BL115 BL_115 bit_cell
X116 VDD VSS WL BL116 BL_116 bit_cell
X117 VDD VSS WL BL117 BL_117 bit_cell
X118 VDD VSS WL BL118 BL_118 bit_cell
X119 VDD VSS WL BL119 BL_119 bit_cell
X120 VDD VSS WL BL120 BL_120 bit_cell
X121 VDD VSS WL BL121 BL_121 bit_cell
X122 VDD VSS WL BL122 BL_122 bit_cell
X123 VDD VSS WL BL123 BL_123 bit_cell
X124 VDD VSS WL BL124 BL_124 bit_cell
X125 VDD VSS WL BL125 BL_125 bit_cell
X126 VDD VSS WL BL126 BL_126 bit_cell
X127 VDD VSS WL BL127 BL_127 bit_cell
.ends bit_arr_128

.subckt dmy_arr_64 VDD VSS WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 WL32 WL33 WL34 WL35 WL36 WL37 WL38 WL39 WL40 WL41 WL42 WL43 WL44 WL45 WL46 WL47 WL48 WL49 WL50 WL51 WL52 WL53 WL54 WL55 WL56 WL57 WL58 WL59 WL60 WL61 WL62 WL63 DBL DBL_
X0 VDD VSS WL0 DBL DBL_ dmy_cell
X1 VDD VSS WL1 DBL DBL_ dmy_cell
X2 VDD VSS WL2 DBL DBL_ dmy_cell
X3 VDD VSS WL3 DBL DBL_ dmy_cell
X4 VDD VSS WL4 DBL DBL_ dmy_cell
X5 VDD VSS WL5 DBL DBL_ dmy_cell
X6 VDD VSS WL6 DBL DBL_ dmy_cell
X7 VDD VSS WL7 DBL DBL_ dmy_cell
X8 VDD VSS WL8 DBL DBL_ dmy_cell
X9 VDD VSS WL9 DBL DBL_ dmy_cell
X10 VDD VSS WL10 DBL DBL_ dmy_cell
X11 VDD VSS WL11 DBL DBL_ dmy_cell
X12 VDD VSS WL12 DBL DBL_ dmy_cell
X13 VDD VSS WL13 DBL DBL_ dmy_cell
X14 VDD VSS WL14 DBL DBL_ dmy_cell
X15 VDD VSS WL15 DBL DBL_ dmy_cell
X16 VDD VSS WL16 DBL DBL_ dmy_cell
X17 VDD VSS WL17 DBL DBL_ dmy_cell
X18 VDD VSS WL18 DBL DBL_ dmy_cell
X19 VDD VSS WL19 DBL DBL_ dmy_cell
X20 VDD VSS WL20 DBL DBL_ dmy_cell
X21 VDD VSS WL21 DBL DBL_ dmy_cell
X22 VDD VSS WL22 DBL DBL_ dmy_cell
X23 VDD VSS WL23 DBL DBL_ dmy_cell
X24 VDD VSS WL24 DBL DBL_ dmy_cell
X25 VDD VSS WL25 DBL DBL_ dmy_cell
X26 VDD VSS WL26 DBL DBL_ dmy_cell
X27 VDD VSS WL27 DBL DBL_ dmy_cell
X28 VDD VSS WL28 DBL DBL_ dmy_cell
X29 VDD VSS WL29 DBL DBL_ dmy_cell
X30 VDD VSS WL30 DBL DBL_ dmy_cell
X31 VDD VSS WL31 DBL DBL_ dmy_cell
X32 VDD VSS WL32 DBL DBL_ dmy_cell
X33 VDD VSS WL33 DBL DBL_ dmy_cell
X34 VDD VSS WL34 DBL DBL_ dmy_cell
X35 VDD VSS WL35 DBL DBL_ dmy_cell
X36 VDD VSS WL36 DBL DBL_ dmy_cell
X37 VDD VSS WL37 DBL DBL_ dmy_cell
X38 VDD VSS WL38 DBL DBL_ dmy_cell
X39 VDD VSS WL39 DBL DBL_ dmy_cell
X40 VDD VSS WL40 DBL DBL_ dmy_cell
X41 VDD VSS WL41 DBL DBL_ dmy_cell
X42 VDD VSS WL42 DBL DBL_ dmy_cell
X43 VDD VSS WL43 DBL DBL_ dmy_cell
X44 VDD VSS WL44 DBL DBL_ dmy_cell
X45 VDD VSS WL45 DBL DBL_ dmy_cell
X46 VDD VSS WL46 DBL DBL_ dmy_cell
X47 VDD VSS WL47 DBL DBL_ dmy_cell
X48 VDD VSS WL48 DBL DBL_ dmy_cell
X49 VDD VSS WL49 DBL DBL_ dmy_cell
X50 VDD VSS WL50 DBL DBL_ dmy_cell
X51 VDD VSS WL51 DBL DBL_ dmy_cell
X52 VDD VSS WL52 DBL DBL_ dmy_cell
X53 VDD VSS WL53 DBL DBL_ dmy_cell
X54 VDD VSS WL54 DBL DBL_ dmy_cell
X55 VDD VSS WL55 DBL DBL_ dmy_cell
X56 VDD VSS WL56 DBL DBL_ dmy_cell
X57 VDD VSS WL57 DBL DBL_ dmy_cell
X58 VDD VSS WL58 DBL DBL_ dmy_cell
X59 VDD VSS WL59 DBL DBL_ dmy_cell
X60 VDD VSS WL60 DBL DBL_ dmy_cell
X61 VDD VSS WL61 DBL DBL_ dmy_cell
X62 VDD VSS WL62 DBL DBL_ dmy_cell
X63 VDD VSS WL63 DBL DBL_ dmy_cell
.ends dmy_arr_64

.subckt se_arr_32 VDD VSS SAEN BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 SB0 SB1 SB2 SB3 SB4 SB5 SB6 SB7 SB8 SB9 SB10 SB11 SB12 SB13 SB14 SB15 SB16 SB17 SB18 SB19 SB20 SB21 SB22 SB23 SB24 SB25 SB26 SB27 SB28 SB29 SB30 SB31
X0 VDD VSS SAEN BL0 BL_0 SB0 se_cell
X1 VDD VSS SAEN BL1 BL_1 SB1 se_cell
X2 VDD VSS SAEN BL2 BL_2 SB2 se_cell
X3 VDD VSS SAEN BL3 BL_3 SB3 se_cell
X4 VDD VSS SAEN BL4 BL_4 SB4 se_cell
X5 VDD VSS SAEN BL5 BL_5 SB5 se_cell
X6 VDD VSS SAEN BL6 BL_6 SB6 se_cell
X7 VDD VSS SAEN BL7 BL_7 SB7 se_cell
X8 VDD VSS SAEN BL8 BL_8 SB8 se_cell
X9 VDD VSS SAEN BL9 BL_9 SB9 se_cell
X10 VDD VSS SAEN BL10 BL_10 SB10 se_cell
X11 VDD VSS SAEN BL11 BL_11 SB11 se_cell
X12 VDD VSS SAEN BL12 BL_12 SB12 se_cell
X13 VDD VSS SAEN BL13 BL_13 SB13 se_cell
X14 VDD VSS SAEN BL14 BL_14 SB14 se_cell
X15 VDD VSS SAEN BL15 BL_15 SB15 se_cell
X16 VDD VSS SAEN BL16 BL_16 SB16 se_cell
X17 VDD VSS SAEN BL17 BL_17 SB17 se_cell
X18 VDD VSS SAEN BL18 BL_18 SB18 se_cell
X19 VDD VSS SAEN BL19 BL_19 SB19 se_cell
X20 VDD VSS SAEN BL20 BL_20 SB20 se_cell
X21 VDD VSS SAEN BL21 BL_21 SB21 se_cell
X22 VDD VSS SAEN BL22 BL_22 SB22 se_cell
X23 VDD VSS SAEN BL23 BL_23 SB23 se_cell
X24 VDD VSS SAEN BL24 BL_24 SB24 se_cell
X25 VDD VSS SAEN BL25 BL_25 SB25 se_cell
X26 VDD VSS SAEN BL26 BL_26 SB26 se_cell
X27 VDD VSS SAEN BL27 BL_27 SB27 se_cell
X28 VDD VSS SAEN BL28 BL_28 SB28 se_cell
X29 VDD VSS SAEN BL29 BL_29 SB29 se_cell
X30 VDD VSS SAEN BL30 BL_30 SB30 se_cell
X31 VDD VSS SAEN BL31 BL_31 SB31 se_cell
.ends se_arr_32

.subckt mat_arr_128 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 WL32 WL33 WL34 WL35 WL36 WL37 WL38 WL39 WL40 WL41 WL42 WL43 WL44 WL45 WL46 WL47 WL48 WL49 WL50 WL51 WL52 WL53 WL54 WL55 WL56 WL57 WL58 WL59 WL60 WL61 WL62 WL63
X0 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL0 bit_arr_128
X1 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL1 bit_arr_128
X2 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL2 bit_arr_128
X3 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL3 bit_arr_128
X4 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL4 bit_arr_128
X5 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL5 bit_arr_128
X6 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL6 bit_arr_128
X7 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL7 bit_arr_128
X8 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL8 bit_arr_128
X9 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL9 bit_arr_128
X10 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL10 bit_arr_128
X11 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL11 bit_arr_128
X12 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL12 bit_arr_128
X13 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL13 bit_arr_128
X14 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL14 bit_arr_128
X15 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL15 bit_arr_128
X16 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL16 bit_arr_128
X17 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL17 bit_arr_128
X18 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL18 bit_arr_128
X19 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL19 bit_arr_128
X20 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL20 bit_arr_128
X21 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL21 bit_arr_128
X22 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL22 bit_arr_128
X23 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL23 bit_arr_128
X24 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL24 bit_arr_128
X25 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL25 bit_arr_128
X26 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL26 bit_arr_128
X27 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL27 bit_arr_128
X28 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL28 bit_arr_128
X29 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL29 bit_arr_128
X30 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL30 bit_arr_128
X31 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL31 bit_arr_128
X32 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL32 bit_arr_128
X33 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL33 bit_arr_128
X34 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL34 bit_arr_128
X35 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL35 bit_arr_128
X36 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL36 bit_arr_128
X37 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL37 bit_arr_128
X38 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL38 bit_arr_128
X39 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL39 bit_arr_128
X40 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL40 bit_arr_128
X41 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL41 bit_arr_128
X42 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL42 bit_arr_128
X43 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL43 bit_arr_128
X44 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL44 bit_arr_128
X45 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL45 bit_arr_128
X46 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL46 bit_arr_128
X47 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL47 bit_arr_128
X48 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL48 bit_arr_128
X49 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL49 bit_arr_128
X50 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL50 bit_arr_128
X51 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL51 bit_arr_128
X52 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL52 bit_arr_128
X53 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL53 bit_arr_128
X54 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL54 bit_arr_128
X55 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL55 bit_arr_128
X56 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL56 bit_arr_128
X57 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL57 bit_arr_128
X58 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL58 bit_arr_128
X59 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL59 bit_arr_128
X60 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL60 bit_arr_128
X61 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL61 bit_arr_128
X62 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL62 bit_arr_128
X63 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL63 bit_arr_128
.ends mat_arr_128

.subckt sram256x32 VDD VSS clk addr0 addr1 addr2 addr3 addr4 addr5 addr6 addr7 din0 din1 din2 din3 din4 din5 din6 din7 din8 din9 din10 din11 din12 din13 din14 din15 din16 din17 din18 din19 din20 din21 din22 din23 din24 din25 din26 din27 din28 din29 din30 din31 Q0 Q1 Q2 Q3 Q4 Q5 Q6 Q7 Q8 Q9 Q10 Q11 Q12 Q13 Q14 Q15 Q16 Q17 Q18 Q19 Q20 Q21 Q22 Q23 Q24 Q25 Q26 Q27 Q28 Q29 Q30 Q31 w_en cs
X0 VDD VSS clk addr0 addr1 addr2 addr3 addr4 addr5 addr6 addr7 w_en A0 A1 A2 A3 A4 A5 A6 A7 write input_reg9
X1 VDD VSS A2 A3 A4 A5 A6 A7 DC0 DC1 DC2 DC3 DC4 DC5 DC6 DC7 DC8 DC9 DC10 DC11 DC12 DC13 DC14 DC15 DC16 DC17 DC18 DC19 DC20 DC21 DC22 DC23 DC24 DC25 DC26 DC27 DC28 DC29 DC30 DC31 DC32 DC33 DC34 DC35 DC36 DC37 DC38 DC39 DC40 DC41 DC42 DC43 DC44 DC45 DC46 DC47 DC48 DC49 DC50 DC51 DC52 DC53 DC54 DC55 DC56 DC57 DC58 DC59 DC60 DC61 DC62 DC63 row_dec64
X2 VDD VSS WLEN DC0 DC1 DC2 DC3 DC4 DC5 DC6 DC7 DC8 DC9 DC10 DC11 DC12 DC13 DC14 DC15 DC16 DC17 DC18 DC19 DC20 DC21 DC22 DC23 DC24 DC25 DC26 DC27 DC28 DC29 DC30 DC31 DC32 DC33 DC34 DC35 DC36 DC37 DC38 DC39 DC40 DC41 DC42 DC43 DC44 DC45 DC46 DC47 DC48 DC49 DC50 DC51 DC52 DC53 DC54 DC55 DC56 DC57 DC58 DC59 DC60 DC61 DC62 DC63 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 WL32 WL33 WL34 WL35 WL36 WL37 WL38 WL39 WL40 WL41 WL42 WL43 WL44 WL45 WL46 WL47 WL48 WL49 WL50 WL51 WL52 WL53 WL54 WL55 WL56 WL57 WL58 WL59 WL60 WL61 WL62 WL63 rd_arr_64
X3 VDD VSS A0 A1 CD0 CD1 CD2 CD3 col_dec4
X4 VDD VSS WLEN CD0 CD1 CD2 CD3 SEL0 SEL1 SEL2 SEL3 rd_arr_4
X5 VDD VSS PCHG WREN SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 DW0 DW_0 DW0 DW_0 DW0 DW_0 DW0 DW_0 DW1 DW_1 DW1 DW_1 DW1 DW_1 DW1 DW_1 DW2 DW_2 DW2 DW_2 DW2 DW_2 DW2 DW_2 DW3 DW_3 DW3 DW_3 DW3 DW_3 DW3 DW_3 DW4 DW_4 DW4 DW_4 DW4 DW_4 DW4 DW_4 DW5 DW_5 DW5 DW_5 DW5 DW_5 DW5 DW_5 DW6 DW_6 DW6 DW_6 DW6 DW_6 DW6 DW_6 DW7 DW_7 DW7 DW_7 DW7 DW_7 DW7 DW_7 DW8 DW_8 DW8 DW_8 DW8 DW_8 DW8 DW_8 DW9 DW_9 DW9 DW_9 DW9 DW_9 DW9 DW_9 DW10 DW_10 DW10 DW_10 DW10 DW_10 DW10 DW_10 DW11 DW_11 DW11 DW_11 DW11 DW_11 DW11 DW_11 DW12 DW_12 DW12 DW_12 DW12 DW_12 DW12 DW_12 DW13 DW_13 DW13 DW_13 DW13 DW_13 DW13 DW_13 DW14 DW_14 DW14 DW_14 DW14 DW_14 DW14 DW_14 DW15 DW_15 DW15 DW_15 DW15 DW_15 DW15 DW_15 DW16 DW_16 DW16 DW_16 DW16 DW_16 DW16 DW_16 DW17 DW_17 DW17 DW_17 DW17 DW_17 DW17 DW_17 DW18 DW_18 DW18 DW_18 DW18 DW_18 DW18 DW_18 DW19 DW_19 DW19 DW_19 DW19 DW_19 DW19 DW_19 DW20 DW_20 DW20 DW_20 DW20 DW_20 DW20 DW_20 DW21 DW_21 DW21 DW_21 DW21 DW_21 DW21 DW_21 DW22 DW_22 DW22 DW_22 DW22 DW_22 DW22 DW_22 DW23 DW_23 DW23 DW_23 DW23 DW_23 DW23 DW_23 DW24 DW_24 DW24 DW_24 DW24 DW_24 DW24 DW_24 DW25 DW_25 DW25 DW_25 DW25 DW_25 DW25 DW_25 DW26 DW_26 DW26 DW_26 DW26 DW_26 DW26 DW_26 DW27 DW_27 DW27 DW_27 DW27 DW_27 DW27 DW_27 DW28 DW_28 DW28 DW_28 DW28 DW_28 DW28 DW_28 DW29 DW_29 DW29 DW_29 DW29 DW_29 DW29 DW_29 DW30 DW_30 DW30 DW_30 DW30 DW_30 DW30 DW_30 DW31 DW_31 DW31 DW_31 DW31 DW_31 DW31 DW_31 DR0 DR_0 DR0 DR_0 DR0 DR_0 DR0 DR_0 DR1 DR_1 DR1 DR_1 DR1 DR_1 DR1 DR_1 DR2 DR_2 DR2 DR_2 DR2 DR_2 DR2 DR_2 DR3 DR_3 DR3 DR_3 DR3 DR_3 DR3 DR_3 DR4 DR_4 DR4 DR_4 DR4 DR_4 DR4 DR_4 DR5 DR_5 DR5 DR_5 DR5 DR_5 DR5 DR_5 DR6 DR_6 DR6 DR_6 DR6 DR_6 DR6 DR_6 DR7 DR_7 DR7 DR_7 DR7 DR_7 DR7 DR_7 DR8 DR_8 DR8 DR_8 DR8 DR_8 DR8 DR_8 DR9 DR_9 DR9 DR_9 DR9 DR_9 DR9 DR_9 DR10 DR_10 DR10 DR_10 DR10 DR_10 DR10 DR_10 DR11 DR_11 DR11 DR_11 DR11 DR_11 DR11 DR_11 DR12 DR_12 DR12 DR_12 DR12 DR_12 DR12 DR_12 DR13 DR_13 DR13 DR_13 DR13 DR_13 DR13 DR_13 DR14 DR_14 DR14 DR_14 DR14 DR_14 DR14 DR_14 DR15 DR_15 DR15 DR_15 DR15 DR_15 DR15 DR_15 DR16 DR_16 DR16 DR_16 DR16 DR_16 DR16 DR_16 DR17 DR_17 DR17 DR_17 DR17 DR_17 DR17 DR_17 DR18 DR_18 DR18 DR_18 DR18 DR_18 DR18 DR_18 DR19 DR_19 DR19 DR_19 DR19 DR_19 DR19 DR_19 DR20 DR_20 DR20 DR_20 DR20 DR_20 DR20 DR_20 DR21 DR_21 DR21 DR_21 DR21 DR_21 DR21 DR_21 DR22 DR_22 DR22 DR_22 DR22 DR_22 DR22 DR_22 DR23 DR_23 DR23 DR_23 DR23 DR_23 DR23 DR_23 DR24 DR_24 DR24 DR_24 DR24 DR_24 DR24 DR_24 DR25 DR_25 DR25 DR_25 DR25 DR_25 DR25 DR_25 DR26 DR_26 DR26 DR_26 DR26 DR_26 DR26 DR_26 DR27 DR_27 DR27 DR_27 DR27 DR_27 DR27 DR_27 DR28 DR_28 DR28 DR_28 DR28 DR_28 DR28 DR_28 DR29 DR_29 DR29 DR_29 DR29 DR_29 DR29 DR_29 DR30 DR_30 DR30 DR_30 DR30 DR_30 DR30 DR_30 DR31 DR_31 DR31 DR_31 DR31 DR_31 DR31 DR_31 dido_arr_128
X6 VDD VSS clk WREN din0 din1 din2 din3 din4 din5 din6 din7 din8 din9 din10 din11 din12 din13 din14 din15 din16 din17 din18 din19 din20 din21 din22 din23 din24 din25 din26 din27 din28 din29 din30 din31 DW0 DW_0 DW1 DW_1 DW2 DW_2 DW3 DW_3 DW4 DW_4 DW5 DW_5 DW6 DW_6 DW7 DW_7 DW8 DW_8 DW9 DW_9 DW10 DW_10 DW11 DW_11 DW12 DW_12 DW13 DW_13 DW14 DW_14 DW15 DW_15 DW16 DW_16 DW17 DW_17 DW18 DW_18 DW19 DW_19 DW20 DW_20 DW21 DW_21 DW22 DW_22 DW23 DW_23 DW24 DW_24 DW25 DW_25 DW26 DW_26 DW27 DW_27 DW28 DW_28 DW29 DW_29 DW30 DW_30 DW31 DW_31 datain_reg32
X7 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 WL32 WL33 WL34 WL35 WL36 WL37 WL38 WL39 WL40 WL41 WL42 WL43 WL44 WL45 WL46 WL47 WL48 WL49 WL50 WL51 WL52 WL53 WL54 WL55 WL56 WL57 WL58 WL59 WL60 WL61 WL62 WL63 mat_arr_128
X8 VDD VSS SAEN DR0 DR_0 DR1 DR_1 DR2 DR_2 DR3 DR_3 DR4 DR_4 DR5 DR_5 DR6 DR_6 DR7 DR_7 DR8 DR_8 DR9 DR_9 DR10 DR_10 DR11 DR_11 DR12 DR_12 DR13 DR_13 DR14 DR_14 DR15 DR_15 DR16 DR_16 DR17 DR_17 DR18 DR_18 DR19 DR_19 DR20 DR_20 DR21 DR_21 DR22 DR_22 DR23 DR_23 DR24 DR_24 DR25 DR_25 DR26 DR_26 DR27 DR_27 DR28 DR_28 DR29 DR_29 DR30 DR_30 DR31 DR_31 Q0 Q1 Q2 Q3 Q4 Q5 Q6 Q7 Q8 Q9 Q10 Q11 Q12 Q13 Q14 Q15 Q16 Q17 Q18 Q19 Q20 Q21 Q22 Q23 Q24 Q25 Q26 Q27 Q28 Q29 Q30 Q31 se_arr_32
X9 VDD VSS clk cs write DBL DBL_ WREN PCHG WLEN SAEN ctrl
X10 VDD VSS WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 WL32 WL33 WL34 WL35 WL36 WL37 WL38 WL39 WL40 WL41 WL42 WL43 WL44 WL45 WL46 WL47 WL48 WL49 WL50 WL51 WL52 WL53 WL54 WL55 WL56 WL57 WL58 WL59 WL60 WL61 WL62 WL63 DBL DBL_ dmy_arr_64
.ends sram256x32

