* SPICE3 file created from sense_amplifier.ext - technology: sky130A

X0 bit_cell_0/a_381_381# bit_cell_0/WL bit_cell_0/BL m9/VSUBS sky130_fd_pr__nfet_01v8 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=0.15
X1 bit_cell_0/a_381_381# bit_cell_0/a_257_458# bit_cell_0/VDD bit_cell_0/VDD sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X2 bit_cell_0/a_257_458# bit_cell_0/a_381_381# bit_cell_0/VDD bit_cell_0/VDD sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.82365 ps=7.43 w=0.42 l=0.15
X3 bit_cell_0/a_381_381# bit_cell_0/a_257_458# m9/VSUBS m9/VSUBS sky130_fd_pr__nfet_01v8 ad=0.232 pd=2.18 as=0.232 ps=2.18 w=0.8 l=0.15
X4 bit_cell_0/a_257_458# bit_cell_0/a_381_381# m9/VSUBS m9/VSUBS sky130_fd_pr__nfet_01v8 ad=0.406 pd=3.96 as=1.05565 ps=9.03 w=0.8 l=0.15
X5 bit_cell_0/BL_ bit_cell_0/WL bit_cell_0/a_257_458# m9/VSUBS sky130_fd_pr__nfet_01v8 ad=0.754 pd=6.36 as=0 ps=0 w=0.6 l=0.15
X6 a_94_n338# a_39_110# m1_136_23# m9/VSUBS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X7 a_286_83# a_182_49# m1_136_23# m9/VSUBS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.365425 ps=3.685 w=0.42 l=0.15
X8 a_94_n338# a_94_n338# bit_cell_0/VDD bit_cell_0/VDD sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X9 a_286_83# a_94_n338# bit_cell_0/VDD bit_cell_0/VDD sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X10 bit_cell_0/BL a_286_83# bit_cell_0/VDD bit_cell_0/VDD sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X11 bit_cell_0/BL a_286_83# m9/VSUBS m9/VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X12 bit_cell_0/BL_ bit_cell_0/BL bit_cell_0/VDD bit_cell_0/VDD sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X13 m1_136_23# a_94_479# m9/VSUBS m9/VSUBS sky130_fd_pr__nfet_01v8 ad=0.2436 pd=2.26 as=0.2436 ps=2.26 w=0.84 l=0.15
X14 bit_cell_0/BL_ bit_cell_0/BL m9/VSUBS m9/VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15
