magic
tech sky130A
magscale 1 2
timestamp 1703060231
<< nwell >>
rect -109 -462 109 462
<< pmos >>
rect -15 -400 15 400
<< pdiff >>
rect -73 388 -15 400
rect -73 -388 -61 388
rect -27 -388 -15 388
rect -73 -400 -15 -388
rect 15 388 73 400
rect 15 -388 27 388
rect 61 -388 73 388
rect 15 -400 73 -388
<< pdiffc >>
rect -61 -388 -27 388
rect 27 -388 61 388
<< poly >>
rect -15 400 15 426
rect -15 -426 15 -400
<< locali >>
rect -61 388 -27 404
rect -61 -404 -27 -388
rect 27 388 61 404
rect 27 -404 61 -388
<< viali >>
rect -61 -388 -27 388
rect 27 -388 61 388
<< metal1 >>
rect -67 388 -21 400
rect -67 -388 -61 388
rect -27 -388 -21 388
rect -67 -400 -21 -388
rect 21 388 67 400
rect 21 -388 27 388
rect 61 -388 67 388
rect 21 -400 67 -388
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
