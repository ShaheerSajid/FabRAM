.title sram_gen
.subckt bit_cell VDD VSS WL BL BL_
X0 Q Q_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X1 Q_ Q VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X2 Q Q_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 Q_ Q VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 Q WL BL VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
X5 Q_ WL BL_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
.ends bit_cell

.subckt dmy_cell VDD VSS WL BL BL_
X0 Q VSS VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X1 Q_ VDD VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X2 Q VSS VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 Q_ VDD VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 Q WL BL VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
X5 Q_ WL BL_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
.ends dmy_cell

.subckt in_reg VDD VSS clk D Q
X0 net3 clk VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X8 net3 clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 net4 net2 net5 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X10 Din net2 net1 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 net55 Q VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X13 net55 Q VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 net2 net3 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X11 net2 net3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X5 Din net3 net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X15 net4 net3 net5 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 Q net5 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X9 Q net5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X6 net11 net4 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X12 net11 net4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X7 net4 net1 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X14 net4 net1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X16 net11 net2 net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X17 net11 net3 net1 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X18 net55 net3 net5 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X19 net55 net2 net5 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X20 D_ D VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X21 D_ D VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X22 Din D_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X23 Din D_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
.ends in_reg

.subckt se_cell VDD VSS SAEN BL BL_ SB
X0 net1 SAEN VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.84
X1 diff1 BL_ net1 net1 sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X2 diff2 BL net1 net1 sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X3 diff1 diff1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 diff2 diff1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X5 diff2_ diff2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X6 diff2_ diff2 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=2
X7 SB_ diff2_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X8 SB_ diff2_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=2
X9 SB_w Q_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X10 Q_ SB_w VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X11 SB_w Q_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X12 Q_ SB_w VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X13 SB_w SAEN SB_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
X14 Q_ SAEN diff2_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
X15 SB SB_w VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X16 SB SB_w VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
.ends se_cell

.subckt not VDD VSS A B
X0 B A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 B A VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends not

.subckt notdel VDD VSS A B
X0 B A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.84
X1 B A VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends notdel

.subckt nand2 VDD VSS A B Y
X0 Y A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 Y B VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 Y B net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X3 net1 A VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends nand2

.subckt nand3 VDD VSS A B C Y
X0 Y A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 Y B VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 Y C VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 Y A net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X4 net1 B net2 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X5 net2 C VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends nand3

.subckt nand4 VDD VSS A B C D Y
X0 Y A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 Y B VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 Y C VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 Y D VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 Y D net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X5 net1 B net2 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X6 net2 C net3 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X7 net3 A VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends nand4

.subckt dec_2to4 VDD VSS A1 A0 Y0 Y1 Y2 Y3
X0 VDD VSS A1 A_1 not
X1 VDD VSS A0 A_0 not
X2 VDD VSS A_1 A_0 Y0_ nand2
X3 VDD VSS A_1 A0 Y1_ nand2
X4 VDD VSS A1 A_0 Y2_ nand2
X5 VDD VSS A1 A0 Y3_ nand2
X6 VDD VSS Y0_ Y0 not
X7 VDD VSS Y1_ Y1 not
X8 VDD VSS Y2_ Y2 not
X9 VDD VSS Y3_ Y3 not
.ends dec_2to4

.subckt dec_3to6 VDD VSS A2 A1 A0 Y0 Y1 Y2 Y3 Y4 Y5
X0 VDD VSS A2 Y4 not
X1 VDD VSS Y4 Y5 not
X2 VDD VSS A1 A0 Y0 Y1 Y2 Y3 dec_2to4
.ends dec_3to6

.subckt row_dec32 VDD VSS A0 A1 A2 A3 A4 DC0 DC1 DC2 DC3 DC4 DC5 DC6 DC7 DC8 DC9 DC10 DC11 DC12 DC13 DC14 DC15 DC16 DC17 DC18 DC19 DC20 DC21 DC22 DC23 DC24 DC25 DC26 DC27 DC28 DC29 DC30 DC31
X0 VDD VSS A1 A0 Y0 Y1 Y2 Y3 dec_2to4
X1 VDD VSS A4 A3 A2 Y4 Y5 Y6 Y7 Y8 Y9 dec_3to6
X2 VDD VSS Y0 Y4 Y8 DC_0 nand3
X3 VDD VSS Y1 Y4 Y8 DC_1 nand3
X4 VDD VSS Y2 Y4 Y8 DC_2 nand3
X5 VDD VSS Y3 Y4 Y8 DC_3 nand3
X6 VDD VSS Y0 Y5 Y8 DC_4 nand3
X7 VDD VSS Y1 Y5 Y8 DC_5 nand3
X8 VDD VSS Y2 Y5 Y8 DC_6 nand3
X9 VDD VSS Y3 Y5 Y8 DC_7 nand3
X10 VDD VSS Y0 Y6 Y8 DC_8 nand3
X11 VDD VSS Y1 Y6 Y8 DC_9 nand3
X12 VDD VSS Y2 Y6 Y8 DC_10 nand3
X13 VDD VSS Y3 Y6 Y8 DC_11 nand3
X14 VDD VSS Y0 Y7 Y8 DC_12 nand3
X15 VDD VSS Y1 Y7 Y8 DC_13 nand3
X16 VDD VSS Y2 Y7 Y8 DC_14 nand3
X17 VDD VSS Y3 Y7 Y8 DC_15 nand3
X18 VDD VSS Y0 Y4 Y9 DC_16 nand3
X19 VDD VSS Y1 Y4 Y9 DC_17 nand3
X20 VDD VSS Y2 Y4 Y9 DC_18 nand3
X21 VDD VSS Y3 Y4 Y9 DC_19 nand3
X22 VDD VSS Y0 Y5 Y9 DC_20 nand3
X23 VDD VSS Y1 Y5 Y9 DC_21 nand3
X24 VDD VSS Y2 Y5 Y9 DC_22 nand3
X25 VDD VSS Y3 Y5 Y9 DC_23 nand3
X26 VDD VSS Y0 Y6 Y9 DC_24 nand3
X27 VDD VSS Y1 Y6 Y9 DC_25 nand3
X28 VDD VSS Y2 Y6 Y9 DC_26 nand3
X29 VDD VSS Y3 Y6 Y9 DC_27 nand3
X30 VDD VSS Y0 Y7 Y9 DC_28 nand3
X31 VDD VSS Y1 Y7 Y9 DC_29 nand3
X32 VDD VSS Y2 Y7 Y9 DC_30 nand3
X33 VDD VSS Y3 Y7 Y9 DC_31 nand3
X34 VDD VSS DC_0 DC0 not
X35 VDD VSS DC_1 DC1 not
X36 VDD VSS DC_2 DC2 not
X37 VDD VSS DC_3 DC3 not
X38 VDD VSS DC_4 DC4 not
X39 VDD VSS DC_5 DC5 not
X40 VDD VSS DC_6 DC6 not
X41 VDD VSS DC_7 DC7 not
X42 VDD VSS DC_8 DC8 not
X43 VDD VSS DC_9 DC9 not
X44 VDD VSS DC_10 DC10 not
X45 VDD VSS DC_11 DC11 not
X46 VDD VSS DC_12 DC12 not
X47 VDD VSS DC_13 DC13 not
X48 VDD VSS DC_14 DC14 not
X49 VDD VSS DC_15 DC15 not
X50 VDD VSS DC_16 DC16 not
X51 VDD VSS DC_17 DC17 not
X52 VDD VSS DC_18 DC18 not
X53 VDD VSS DC_19 DC19 not
X54 VDD VSS DC_20 DC20 not
X55 VDD VSS DC_21 DC21 not
X56 VDD VSS DC_22 DC22 not
X57 VDD VSS DC_23 DC23 not
X58 VDD VSS DC_24 DC24 not
X59 VDD VSS DC_25 DC25 not
X60 VDD VSS DC_26 DC26 not
X61 VDD VSS DC_27 DC27 not
X62 VDD VSS DC_28 DC28 not
X63 VDD VSS DC_29 DC29 not
X64 VDD VSS DC_30 DC30 not
X65 VDD VSS DC_31 DC31 not
.ends row_dec32

.subckt row_driver VDD VSS WLEN A B
X0 VDD VSS A WLEN net1 nand2
X1 B net1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X2 B net1 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
.ends row_driver

.subckt rd_arr_32 VDD VSS WLEN DC0 DC1 DC2 DC3 DC4 DC5 DC6 DC7 DC8 DC9 DC10 DC11 DC12 DC13 DC14 DC15 DC16 DC17 DC18 DC19 DC20 DC21 DC22 DC23 DC24 DC25 DC26 DC27 DC28 DC29 DC30 DC31 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31
X0 VDD VSS WLEN DC0 WL0 row_driver
X1 VDD VSS WLEN DC1 WL1 row_driver
X2 VDD VSS WLEN DC2 WL2 row_driver
X3 VDD VSS WLEN DC3 WL3 row_driver
X4 VDD VSS WLEN DC4 WL4 row_driver
X5 VDD VSS WLEN DC5 WL5 row_driver
X6 VDD VSS WLEN DC6 WL6 row_driver
X7 VDD VSS WLEN DC7 WL7 row_driver
X8 VDD VSS WLEN DC8 WL8 row_driver
X9 VDD VSS WLEN DC9 WL9 row_driver
X10 VDD VSS WLEN DC10 WL10 row_driver
X11 VDD VSS WLEN DC11 WL11 row_driver
X12 VDD VSS WLEN DC12 WL12 row_driver
X13 VDD VSS WLEN DC13 WL13 row_driver
X14 VDD VSS WLEN DC14 WL14 row_driver
X15 VDD VSS WLEN DC15 WL15 row_driver
X16 VDD VSS WLEN DC16 WL16 row_driver
X17 VDD VSS WLEN DC17 WL17 row_driver
X18 VDD VSS WLEN DC18 WL18 row_driver
X19 VDD VSS WLEN DC19 WL19 row_driver
X20 VDD VSS WLEN DC20 WL20 row_driver
X21 VDD VSS WLEN DC21 WL21 row_driver
X22 VDD VSS WLEN DC22 WL22 row_driver
X23 VDD VSS WLEN DC23 WL23 row_driver
X24 VDD VSS WLEN DC24 WL24 row_driver
X25 VDD VSS WLEN DC25 WL25 row_driver
X26 VDD VSS WLEN DC26 WL26 row_driver
X27 VDD VSS WLEN DC27 WL27 row_driver
X28 VDD VSS WLEN DC28 WL28 row_driver
X29 VDD VSS WLEN DC29 WL29 row_driver
X30 VDD VSS WLEN DC30 WL30 row_driver
X31 VDD VSS WLEN DC31 WL31 row_driver
.ends rd_arr_32

.subckt rd_arr_4 VDD VSS WLEN DC0 DC1 DC2 DC3 WL0 WL1 WL2 WL3
X0 VDD VSS WLEN DC0 WL0 row_driver
X1 VDD VSS WLEN DC1 WL1 row_driver
X2 VDD VSS WLEN DC2 WL2 row_driver
X3 VDD VSS WLEN DC3 WL3 row_driver
.ends rd_arr_4

.subckt col_dec4 VDD VSS A0 A1 DC0 DC1 DC2 DC3
X0 VDD VSS A1 A0 Y0 Y1 Y2 Y3 dec_2to4
X1 VDD VSS Y0 DC0 not
X2 VDD VSS Y1 DC1 not
X3 VDD VSS Y2 DC2 not
X4 VDD VSS Y3 DC3 not
.ends col_dec4

.subckt dido VDD VSS PCHG WREN SEL BL BL_ DW DW_ DR DR_
X0 BL_ net6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 BL net6 BL_ VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 BL net6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 net6 net5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 net6 net5 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X5 net5 PCHG VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X6 net5 PCHG VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X7 BL_ net4 DR_ VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X8 DR net4 BL VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X9 net4 SEL VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X10 BL net2 DW VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X11 DW_ net2 BL_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X12 net4 SEL VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X13 net3 net4 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X14 net3 net4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X15 VDD VSS net3 WREN net1 nand2
X16 VDD VSS net1 net2 not
.ends dido

.subckt dido_arr_512 VDD VSS PCHG WREN SEL0 SEL1 SEL2 SEL3 SEL4 SEL5 SEL6 SEL7 SEL8 SEL9 SEL10 SEL11 SEL12 SEL13 SEL14 SEL15 SEL16 SEL17 SEL18 SEL19 SEL20 SEL21 SEL22 SEL23 SEL24 SEL25 SEL26 SEL27 SEL28 SEL29 SEL30 SEL31 SEL32 SEL33 SEL34 SEL35 SEL36 SEL37 SEL38 SEL39 SEL40 SEL41 SEL42 SEL43 SEL44 SEL45 SEL46 SEL47 SEL48 SEL49 SEL50 SEL51 SEL52 SEL53 SEL54 SEL55 SEL56 SEL57 SEL58 SEL59 SEL60 SEL61 SEL62 SEL63 SEL64 SEL65 SEL66 SEL67 SEL68 SEL69 SEL70 SEL71 SEL72 SEL73 SEL74 SEL75 SEL76 SEL77 SEL78 SEL79 SEL80 SEL81 SEL82 SEL83 SEL84 SEL85 SEL86 SEL87 SEL88 SEL89 SEL90 SEL91 SEL92 SEL93 SEL94 SEL95 SEL96 SEL97 SEL98 SEL99 SEL100 SEL101 SEL102 SEL103 SEL104 SEL105 SEL106 SEL107 SEL108 SEL109 SEL110 SEL111 SEL112 SEL113 SEL114 SEL115 SEL116 SEL117 SEL118 SEL119 SEL120 SEL121 SEL122 SEL123 SEL124 SEL125 SEL126 SEL127 SEL128 SEL129 SEL130 SEL131 SEL132 SEL133 SEL134 SEL135 SEL136 SEL137 SEL138 SEL139 SEL140 SEL141 SEL142 SEL143 SEL144 SEL145 SEL146 SEL147 SEL148 SEL149 SEL150 SEL151 SEL152 SEL153 SEL154 SEL155 SEL156 SEL157 SEL158 SEL159 SEL160 SEL161 SEL162 SEL163 SEL164 SEL165 SEL166 SEL167 SEL168 SEL169 SEL170 SEL171 SEL172 SEL173 SEL174 SEL175 SEL176 SEL177 SEL178 SEL179 SEL180 SEL181 SEL182 SEL183 SEL184 SEL185 SEL186 SEL187 SEL188 SEL189 SEL190 SEL191 SEL192 SEL193 SEL194 SEL195 SEL196 SEL197 SEL198 SEL199 SEL200 SEL201 SEL202 SEL203 SEL204 SEL205 SEL206 SEL207 SEL208 SEL209 SEL210 SEL211 SEL212 SEL213 SEL214 SEL215 SEL216 SEL217 SEL218 SEL219 SEL220 SEL221 SEL222 SEL223 SEL224 SEL225 SEL226 SEL227 SEL228 SEL229 SEL230 SEL231 SEL232 SEL233 SEL234 SEL235 SEL236 SEL237 SEL238 SEL239 SEL240 SEL241 SEL242 SEL243 SEL244 SEL245 SEL246 SEL247 SEL248 SEL249 SEL250 SEL251 SEL252 SEL253 SEL254 SEL255 SEL256 SEL257 SEL258 SEL259 SEL260 SEL261 SEL262 SEL263 SEL264 SEL265 SEL266 SEL267 SEL268 SEL269 SEL270 SEL271 SEL272 SEL273 SEL274 SEL275 SEL276 SEL277 SEL278 SEL279 SEL280 SEL281 SEL282 SEL283 SEL284 SEL285 SEL286 SEL287 SEL288 SEL289 SEL290 SEL291 SEL292 SEL293 SEL294 SEL295 SEL296 SEL297 SEL298 SEL299 SEL300 SEL301 SEL302 SEL303 SEL304 SEL305 SEL306 SEL307 SEL308 SEL309 SEL310 SEL311 SEL312 SEL313 SEL314 SEL315 SEL316 SEL317 SEL318 SEL319 SEL320 SEL321 SEL322 SEL323 SEL324 SEL325 SEL326 SEL327 SEL328 SEL329 SEL330 SEL331 SEL332 SEL333 SEL334 SEL335 SEL336 SEL337 SEL338 SEL339 SEL340 SEL341 SEL342 SEL343 SEL344 SEL345 SEL346 SEL347 SEL348 SEL349 SEL350 SEL351 SEL352 SEL353 SEL354 SEL355 SEL356 SEL357 SEL358 SEL359 SEL360 SEL361 SEL362 SEL363 SEL364 SEL365 SEL366 SEL367 SEL368 SEL369 SEL370 SEL371 SEL372 SEL373 SEL374 SEL375 SEL376 SEL377 SEL378 SEL379 SEL380 SEL381 SEL382 SEL383 SEL384 SEL385 SEL386 SEL387 SEL388 SEL389 SEL390 SEL391 SEL392 SEL393 SEL394 SEL395 SEL396 SEL397 SEL398 SEL399 SEL400 SEL401 SEL402 SEL403 SEL404 SEL405 SEL406 SEL407 SEL408 SEL409 SEL410 SEL411 SEL412 SEL413 SEL414 SEL415 SEL416 SEL417 SEL418 SEL419 SEL420 SEL421 SEL422 SEL423 SEL424 SEL425 SEL426 SEL427 SEL428 SEL429 SEL430 SEL431 SEL432 SEL433 SEL434 SEL435 SEL436 SEL437 SEL438 SEL439 SEL440 SEL441 SEL442 SEL443 SEL444 SEL445 SEL446 SEL447 SEL448 SEL449 SEL450 SEL451 SEL452 SEL453 SEL454 SEL455 SEL456 SEL457 SEL458 SEL459 SEL460 SEL461 SEL462 SEL463 SEL464 SEL465 SEL466 SEL467 SEL468 SEL469 SEL470 SEL471 SEL472 SEL473 SEL474 SEL475 SEL476 SEL477 SEL478 SEL479 SEL480 SEL481 SEL482 SEL483 SEL484 SEL485 SEL486 SEL487 SEL488 SEL489 SEL490 SEL491 SEL492 SEL493 SEL494 SEL495 SEL496 SEL497 SEL498 SEL499 SEL500 SEL501 SEL502 SEL503 SEL504 SEL505 SEL506 SEL507 SEL508 SEL509 SEL510 SEL511 BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 DW0 DW_0 DW1 DW_1 DW2 DW_2 DW3 DW_3 DW4 DW_4 DW5 DW_5 DW6 DW_6 DW7 DW_7 DW8 DW_8 DW9 DW_9 DW10 DW_10 DW11 DW_11 DW12 DW_12 DW13 DW_13 DW14 DW_14 DW15 DW_15 DW16 DW_16 DW17 DW_17 DW18 DW_18 DW19 DW_19 DW20 DW_20 DW21 DW_21 DW22 DW_22 DW23 DW_23 DW24 DW_24 DW25 DW_25 DW26 DW_26 DW27 DW_27 DW28 DW_28 DW29 DW_29 DW30 DW_30 DW31 DW_31 DW32 DW_32 DW33 DW_33 DW34 DW_34 DW35 DW_35 DW36 DW_36 DW37 DW_37 DW38 DW_38 DW39 DW_39 DW40 DW_40 DW41 DW_41 DW42 DW_42 DW43 DW_43 DW44 DW_44 DW45 DW_45 DW46 DW_46 DW47 DW_47 DW48 DW_48 DW49 DW_49 DW50 DW_50 DW51 DW_51 DW52 DW_52 DW53 DW_53 DW54 DW_54 DW55 DW_55 DW56 DW_56 DW57 DW_57 DW58 DW_58 DW59 DW_59 DW60 DW_60 DW61 DW_61 DW62 DW_62 DW63 DW_63 DW64 DW_64 DW65 DW_65 DW66 DW_66 DW67 DW_67 DW68 DW_68 DW69 DW_69 DW70 DW_70 DW71 DW_71 DW72 DW_72 DW73 DW_73 DW74 DW_74 DW75 DW_75 DW76 DW_76 DW77 DW_77 DW78 DW_78 DW79 DW_79 DW80 DW_80 DW81 DW_81 DW82 DW_82 DW83 DW_83 DW84 DW_84 DW85 DW_85 DW86 DW_86 DW87 DW_87 DW88 DW_88 DW89 DW_89 DW90 DW_90 DW91 DW_91 DW92 DW_92 DW93 DW_93 DW94 DW_94 DW95 DW_95 DW96 DW_96 DW97 DW_97 DW98 DW_98 DW99 DW_99 DW100 DW_100 DW101 DW_101 DW102 DW_102 DW103 DW_103 DW104 DW_104 DW105 DW_105 DW106 DW_106 DW107 DW_107 DW108 DW_108 DW109 DW_109 DW110 DW_110 DW111 DW_111 DW112 DW_112 DW113 DW_113 DW114 DW_114 DW115 DW_115 DW116 DW_116 DW117 DW_117 DW118 DW_118 DW119 DW_119 DW120 DW_120 DW121 DW_121 DW122 DW_122 DW123 DW_123 DW124 DW_124 DW125 DW_125 DW126 DW_126 DW127 DW_127 DW128 DW_128 DW129 DW_129 DW130 DW_130 DW131 DW_131 DW132 DW_132 DW133 DW_133 DW134 DW_134 DW135 DW_135 DW136 DW_136 DW137 DW_137 DW138 DW_138 DW139 DW_139 DW140 DW_140 DW141 DW_141 DW142 DW_142 DW143 DW_143 DW144 DW_144 DW145 DW_145 DW146 DW_146 DW147 DW_147 DW148 DW_148 DW149 DW_149 DW150 DW_150 DW151 DW_151 DW152 DW_152 DW153 DW_153 DW154 DW_154 DW155 DW_155 DW156 DW_156 DW157 DW_157 DW158 DW_158 DW159 DW_159 DW160 DW_160 DW161 DW_161 DW162 DW_162 DW163 DW_163 DW164 DW_164 DW165 DW_165 DW166 DW_166 DW167 DW_167 DW168 DW_168 DW169 DW_169 DW170 DW_170 DW171 DW_171 DW172 DW_172 DW173 DW_173 DW174 DW_174 DW175 DW_175 DW176 DW_176 DW177 DW_177 DW178 DW_178 DW179 DW_179 DW180 DW_180 DW181 DW_181 DW182 DW_182 DW183 DW_183 DW184 DW_184 DW185 DW_185 DW186 DW_186 DW187 DW_187 DW188 DW_188 DW189 DW_189 DW190 DW_190 DW191 DW_191 DW192 DW_192 DW193 DW_193 DW194 DW_194 DW195 DW_195 DW196 DW_196 DW197 DW_197 DW198 DW_198 DW199 DW_199 DW200 DW_200 DW201 DW_201 DW202 DW_202 DW203 DW_203 DW204 DW_204 DW205 DW_205 DW206 DW_206 DW207 DW_207 DW208 DW_208 DW209 DW_209 DW210 DW_210 DW211 DW_211 DW212 DW_212 DW213 DW_213 DW214 DW_214 DW215 DW_215 DW216 DW_216 DW217 DW_217 DW218 DW_218 DW219 DW_219 DW220 DW_220 DW221 DW_221 DW222 DW_222 DW223 DW_223 DW224 DW_224 DW225 DW_225 DW226 DW_226 DW227 DW_227 DW228 DW_228 DW229 DW_229 DW230 DW_230 DW231 DW_231 DW232 DW_232 DW233 DW_233 DW234 DW_234 DW235 DW_235 DW236 DW_236 DW237 DW_237 DW238 DW_238 DW239 DW_239 DW240 DW_240 DW241 DW_241 DW242 DW_242 DW243 DW_243 DW244 DW_244 DW245 DW_245 DW246 DW_246 DW247 DW_247 DW248 DW_248 DW249 DW_249 DW250 DW_250 DW251 DW_251 DW252 DW_252 DW253 DW_253 DW254 DW_254 DW255 DW_255 DW256 DW_256 DW257 DW_257 DW258 DW_258 DW259 DW_259 DW260 DW_260 DW261 DW_261 DW262 DW_262 DW263 DW_263 DW264 DW_264 DW265 DW_265 DW266 DW_266 DW267 DW_267 DW268 DW_268 DW269 DW_269 DW270 DW_270 DW271 DW_271 DW272 DW_272 DW273 DW_273 DW274 DW_274 DW275 DW_275 DW276 DW_276 DW277 DW_277 DW278 DW_278 DW279 DW_279 DW280 DW_280 DW281 DW_281 DW282 DW_282 DW283 DW_283 DW284 DW_284 DW285 DW_285 DW286 DW_286 DW287 DW_287 DW288 DW_288 DW289 DW_289 DW290 DW_290 DW291 DW_291 DW292 DW_292 DW293 DW_293 DW294 DW_294 DW295 DW_295 DW296 DW_296 DW297 DW_297 DW298 DW_298 DW299 DW_299 DW300 DW_300 DW301 DW_301 DW302 DW_302 DW303 DW_303 DW304 DW_304 DW305 DW_305 DW306 DW_306 DW307 DW_307 DW308 DW_308 DW309 DW_309 DW310 DW_310 DW311 DW_311 DW312 DW_312 DW313 DW_313 DW314 DW_314 DW315 DW_315 DW316 DW_316 DW317 DW_317 DW318 DW_318 DW319 DW_319 DW320 DW_320 DW321 DW_321 DW322 DW_322 DW323 DW_323 DW324 DW_324 DW325 DW_325 DW326 DW_326 DW327 DW_327 DW328 DW_328 DW329 DW_329 DW330 DW_330 DW331 DW_331 DW332 DW_332 DW333 DW_333 DW334 DW_334 DW335 DW_335 DW336 DW_336 DW337 DW_337 DW338 DW_338 DW339 DW_339 DW340 DW_340 DW341 DW_341 DW342 DW_342 DW343 DW_343 DW344 DW_344 DW345 DW_345 DW346 DW_346 DW347 DW_347 DW348 DW_348 DW349 DW_349 DW350 DW_350 DW351 DW_351 DW352 DW_352 DW353 DW_353 DW354 DW_354 DW355 DW_355 DW356 DW_356 DW357 DW_357 DW358 DW_358 DW359 DW_359 DW360 DW_360 DW361 DW_361 DW362 DW_362 DW363 DW_363 DW364 DW_364 DW365 DW_365 DW366 DW_366 DW367 DW_367 DW368 DW_368 DW369 DW_369 DW370 DW_370 DW371 DW_371 DW372 DW_372 DW373 DW_373 DW374 DW_374 DW375 DW_375 DW376 DW_376 DW377 DW_377 DW378 DW_378 DW379 DW_379 DW380 DW_380 DW381 DW_381 DW382 DW_382 DW383 DW_383 DW384 DW_384 DW385 DW_385 DW386 DW_386 DW387 DW_387 DW388 DW_388 DW389 DW_389 DW390 DW_390 DW391 DW_391 DW392 DW_392 DW393 DW_393 DW394 DW_394 DW395 DW_395 DW396 DW_396 DW397 DW_397 DW398 DW_398 DW399 DW_399 DW400 DW_400 DW401 DW_401 DW402 DW_402 DW403 DW_403 DW404 DW_404 DW405 DW_405 DW406 DW_406 DW407 DW_407 DW408 DW_408 DW409 DW_409 DW410 DW_410 DW411 DW_411 DW412 DW_412 DW413 DW_413 DW414 DW_414 DW415 DW_415 DW416 DW_416 DW417 DW_417 DW418 DW_418 DW419 DW_419 DW420 DW_420 DW421 DW_421 DW422 DW_422 DW423 DW_423 DW424 DW_424 DW425 DW_425 DW426 DW_426 DW427 DW_427 DW428 DW_428 DW429 DW_429 DW430 DW_430 DW431 DW_431 DW432 DW_432 DW433 DW_433 DW434 DW_434 DW435 DW_435 DW436 DW_436 DW437 DW_437 DW438 DW_438 DW439 DW_439 DW440 DW_440 DW441 DW_441 DW442 DW_442 DW443 DW_443 DW444 DW_444 DW445 DW_445 DW446 DW_446 DW447 DW_447 DW448 DW_448 DW449 DW_449 DW450 DW_450 DW451 DW_451 DW452 DW_452 DW453 DW_453 DW454 DW_454 DW455 DW_455 DW456 DW_456 DW457 DW_457 DW458 DW_458 DW459 DW_459 DW460 DW_460 DW461 DW_461 DW462 DW_462 DW463 DW_463 DW464 DW_464 DW465 DW_465 DW466 DW_466 DW467 DW_467 DW468 DW_468 DW469 DW_469 DW470 DW_470 DW471 DW_471 DW472 DW_472 DW473 DW_473 DW474 DW_474 DW475 DW_475 DW476 DW_476 DW477 DW_477 DW478 DW_478 DW479 DW_479 DW480 DW_480 DW481 DW_481 DW482 DW_482 DW483 DW_483 DW484 DW_484 DW485 DW_485 DW486 DW_486 DW487 DW_487 DW488 DW_488 DW489 DW_489 DW490 DW_490 DW491 DW_491 DW492 DW_492 DW493 DW_493 DW494 DW_494 DW495 DW_495 DW496 DW_496 DW497 DW_497 DW498 DW_498 DW499 DW_499 DW500 DW_500 DW501 DW_501 DW502 DW_502 DW503 DW_503 DW504 DW_504 DW505 DW_505 DW506 DW_506 DW507 DW_507 DW508 DW_508 DW509 DW_509 DW510 DW_510 DW511 DW_511 DR0 DR_0 DR1 DR_1 DR2 DR_2 DR3 DR_3 DR4 DR_4 DR5 DR_5 DR6 DR_6 DR7 DR_7 DR8 DR_8 DR9 DR_9 DR10 DR_10 DR11 DR_11 DR12 DR_12 DR13 DR_13 DR14 DR_14 DR15 DR_15 DR16 DR_16 DR17 DR_17 DR18 DR_18 DR19 DR_19 DR20 DR_20 DR21 DR_21 DR22 DR_22 DR23 DR_23 DR24 DR_24 DR25 DR_25 DR26 DR_26 DR27 DR_27 DR28 DR_28 DR29 DR_29 DR30 DR_30 DR31 DR_31 DR32 DR_32 DR33 DR_33 DR34 DR_34 DR35 DR_35 DR36 DR_36 DR37 DR_37 DR38 DR_38 DR39 DR_39 DR40 DR_40 DR41 DR_41 DR42 DR_42 DR43 DR_43 DR44 DR_44 DR45 DR_45 DR46 DR_46 DR47 DR_47 DR48 DR_48 DR49 DR_49 DR50 DR_50 DR51 DR_51 DR52 DR_52 DR53 DR_53 DR54 DR_54 DR55 DR_55 DR56 DR_56 DR57 DR_57 DR58 DR_58 DR59 DR_59 DR60 DR_60 DR61 DR_61 DR62 DR_62 DR63 DR_63 DR64 DR_64 DR65 DR_65 DR66 DR_66 DR67 DR_67 DR68 DR_68 DR69 DR_69 DR70 DR_70 DR71 DR_71 DR72 DR_72 DR73 DR_73 DR74 DR_74 DR75 DR_75 DR76 DR_76 DR77 DR_77 DR78 DR_78 DR79 DR_79 DR80 DR_80 DR81 DR_81 DR82 DR_82 DR83 DR_83 DR84 DR_84 DR85 DR_85 DR86 DR_86 DR87 DR_87 DR88 DR_88 DR89 DR_89 DR90 DR_90 DR91 DR_91 DR92 DR_92 DR93 DR_93 DR94 DR_94 DR95 DR_95 DR96 DR_96 DR97 DR_97 DR98 DR_98 DR99 DR_99 DR100 DR_100 DR101 DR_101 DR102 DR_102 DR103 DR_103 DR104 DR_104 DR105 DR_105 DR106 DR_106 DR107 DR_107 DR108 DR_108 DR109 DR_109 DR110 DR_110 DR111 DR_111 DR112 DR_112 DR113 DR_113 DR114 DR_114 DR115 DR_115 DR116 DR_116 DR117 DR_117 DR118 DR_118 DR119 DR_119 DR120 DR_120 DR121 DR_121 DR122 DR_122 DR123 DR_123 DR124 DR_124 DR125 DR_125 DR126 DR_126 DR127 DR_127 DR128 DR_128 DR129 DR_129 DR130 DR_130 DR131 DR_131 DR132 DR_132 DR133 DR_133 DR134 DR_134 DR135 DR_135 DR136 DR_136 DR137 DR_137 DR138 DR_138 DR139 DR_139 DR140 DR_140 DR141 DR_141 DR142 DR_142 DR143 DR_143 DR144 DR_144 DR145 DR_145 DR146 DR_146 DR147 DR_147 DR148 DR_148 DR149 DR_149 DR150 DR_150 DR151 DR_151 DR152 DR_152 DR153 DR_153 DR154 DR_154 DR155 DR_155 DR156 DR_156 DR157 DR_157 DR158 DR_158 DR159 DR_159 DR160 DR_160 DR161 DR_161 DR162 DR_162 DR163 DR_163 DR164 DR_164 DR165 DR_165 DR166 DR_166 DR167 DR_167 DR168 DR_168 DR169 DR_169 DR170 DR_170 DR171 DR_171 DR172 DR_172 DR173 DR_173 DR174 DR_174 DR175 DR_175 DR176 DR_176 DR177 DR_177 DR178 DR_178 DR179 DR_179 DR180 DR_180 DR181 DR_181 DR182 DR_182 DR183 DR_183 DR184 DR_184 DR185 DR_185 DR186 DR_186 DR187 DR_187 DR188 DR_188 DR189 DR_189 DR190 DR_190 DR191 DR_191 DR192 DR_192 DR193 DR_193 DR194 DR_194 DR195 DR_195 DR196 DR_196 DR197 DR_197 DR198 DR_198 DR199 DR_199 DR200 DR_200 DR201 DR_201 DR202 DR_202 DR203 DR_203 DR204 DR_204 DR205 DR_205 DR206 DR_206 DR207 DR_207 DR208 DR_208 DR209 DR_209 DR210 DR_210 DR211 DR_211 DR212 DR_212 DR213 DR_213 DR214 DR_214 DR215 DR_215 DR216 DR_216 DR217 DR_217 DR218 DR_218 DR219 DR_219 DR220 DR_220 DR221 DR_221 DR222 DR_222 DR223 DR_223 DR224 DR_224 DR225 DR_225 DR226 DR_226 DR227 DR_227 DR228 DR_228 DR229 DR_229 DR230 DR_230 DR231 DR_231 DR232 DR_232 DR233 DR_233 DR234 DR_234 DR235 DR_235 DR236 DR_236 DR237 DR_237 DR238 DR_238 DR239 DR_239 DR240 DR_240 DR241 DR_241 DR242 DR_242 DR243 DR_243 DR244 DR_244 DR245 DR_245 DR246 DR_246 DR247 DR_247 DR248 DR_248 DR249 DR_249 DR250 DR_250 DR251 DR_251 DR252 DR_252 DR253 DR_253 DR254 DR_254 DR255 DR_255 DR256 DR_256 DR257 DR_257 DR258 DR_258 DR259 DR_259 DR260 DR_260 DR261 DR_261 DR262 DR_262 DR263 DR_263 DR264 DR_264 DR265 DR_265 DR266 DR_266 DR267 DR_267 DR268 DR_268 DR269 DR_269 DR270 DR_270 DR271 DR_271 DR272 DR_272 DR273 DR_273 DR274 DR_274 DR275 DR_275 DR276 DR_276 DR277 DR_277 DR278 DR_278 DR279 DR_279 DR280 DR_280 DR281 DR_281 DR282 DR_282 DR283 DR_283 DR284 DR_284 DR285 DR_285 DR286 DR_286 DR287 DR_287 DR288 DR_288 DR289 DR_289 DR290 DR_290 DR291 DR_291 DR292 DR_292 DR293 DR_293 DR294 DR_294 DR295 DR_295 DR296 DR_296 DR297 DR_297 DR298 DR_298 DR299 DR_299 DR300 DR_300 DR301 DR_301 DR302 DR_302 DR303 DR_303 DR304 DR_304 DR305 DR_305 DR306 DR_306 DR307 DR_307 DR308 DR_308 DR309 DR_309 DR310 DR_310 DR311 DR_311 DR312 DR_312 DR313 DR_313 DR314 DR_314 DR315 DR_315 DR316 DR_316 DR317 DR_317 DR318 DR_318 DR319 DR_319 DR320 DR_320 DR321 DR_321 DR322 DR_322 DR323 DR_323 DR324 DR_324 DR325 DR_325 DR326 DR_326 DR327 DR_327 DR328 DR_328 DR329 DR_329 DR330 DR_330 DR331 DR_331 DR332 DR_332 DR333 DR_333 DR334 DR_334 DR335 DR_335 DR336 DR_336 DR337 DR_337 DR338 DR_338 DR339 DR_339 DR340 DR_340 DR341 DR_341 DR342 DR_342 DR343 DR_343 DR344 DR_344 DR345 DR_345 DR346 DR_346 DR347 DR_347 DR348 DR_348 DR349 DR_349 DR350 DR_350 DR351 DR_351 DR352 DR_352 DR353 DR_353 DR354 DR_354 DR355 DR_355 DR356 DR_356 DR357 DR_357 DR358 DR_358 DR359 DR_359 DR360 DR_360 DR361 DR_361 DR362 DR_362 DR363 DR_363 DR364 DR_364 DR365 DR_365 DR366 DR_366 DR367 DR_367 DR368 DR_368 DR369 DR_369 DR370 DR_370 DR371 DR_371 DR372 DR_372 DR373 DR_373 DR374 DR_374 DR375 DR_375 DR376 DR_376 DR377 DR_377 DR378 DR_378 DR379 DR_379 DR380 DR_380 DR381 DR_381 DR382 DR_382 DR383 DR_383 DR384 DR_384 DR385 DR_385 DR386 DR_386 DR387 DR_387 DR388 DR_388 DR389 DR_389 DR390 DR_390 DR391 DR_391 DR392 DR_392 DR393 DR_393 DR394 DR_394 DR395 DR_395 DR396 DR_396 DR397 DR_397 DR398 DR_398 DR399 DR_399 DR400 DR_400 DR401 DR_401 DR402 DR_402 DR403 DR_403 DR404 DR_404 DR405 DR_405 DR406 DR_406 DR407 DR_407 DR408 DR_408 DR409 DR_409 DR410 DR_410 DR411 DR_411 DR412 DR_412 DR413 DR_413 DR414 DR_414 DR415 DR_415 DR416 DR_416 DR417 DR_417 DR418 DR_418 DR419 DR_419 DR420 DR_420 DR421 DR_421 DR422 DR_422 DR423 DR_423 DR424 DR_424 DR425 DR_425 DR426 DR_426 DR427 DR_427 DR428 DR_428 DR429 DR_429 DR430 DR_430 DR431 DR_431 DR432 DR_432 DR433 DR_433 DR434 DR_434 DR435 DR_435 DR436 DR_436 DR437 DR_437 DR438 DR_438 DR439 DR_439 DR440 DR_440 DR441 DR_441 DR442 DR_442 DR443 DR_443 DR444 DR_444 DR445 DR_445 DR446 DR_446 DR447 DR_447 DR448 DR_448 DR449 DR_449 DR450 DR_450 DR451 DR_451 DR452 DR_452 DR453 DR_453 DR454 DR_454 DR455 DR_455 DR456 DR_456 DR457 DR_457 DR458 DR_458 DR459 DR_459 DR460 DR_460 DR461 DR_461 DR462 DR_462 DR463 DR_463 DR464 DR_464 DR465 DR_465 DR466 DR_466 DR467 DR_467 DR468 DR_468 DR469 DR_469 DR470 DR_470 DR471 DR_471 DR472 DR_472 DR473 DR_473 DR474 DR_474 DR475 DR_475 DR476 DR_476 DR477 DR_477 DR478 DR_478 DR479 DR_479 DR480 DR_480 DR481 DR_481 DR482 DR_482 DR483 DR_483 DR484 DR_484 DR485 DR_485 DR486 DR_486 DR487 DR_487 DR488 DR_488 DR489 DR_489 DR490 DR_490 DR491 DR_491 DR492 DR_492 DR493 DR_493 DR494 DR_494 DR495 DR_495 DR496 DR_496 DR497 DR_497 DR498 DR_498 DR499 DR_499 DR500 DR_500 DR501 DR_501 DR502 DR_502 DR503 DR_503 DR504 DR_504 DR505 DR_505 DR506 DR_506 DR507 DR_507 DR508 DR_508 DR509 DR_509 DR510 DR_510 DR511 DR_511
X0 VDD VSS PCHG WREN SEL0 BL0 BL_0 DW0 DW_0 DR0 DR_0 dido
X1 VDD VSS PCHG WREN SEL1 BL1 BL_1 DW1 DW_1 DR1 DR_1 dido
X2 VDD VSS PCHG WREN SEL2 BL2 BL_2 DW2 DW_2 DR2 DR_2 dido
X3 VDD VSS PCHG WREN SEL3 BL3 BL_3 DW3 DW_3 DR3 DR_3 dido
X4 VDD VSS PCHG WREN SEL4 BL4 BL_4 DW4 DW_4 DR4 DR_4 dido
X5 VDD VSS PCHG WREN SEL5 BL5 BL_5 DW5 DW_5 DR5 DR_5 dido
X6 VDD VSS PCHG WREN SEL6 BL6 BL_6 DW6 DW_6 DR6 DR_6 dido
X7 VDD VSS PCHG WREN SEL7 BL7 BL_7 DW7 DW_7 DR7 DR_7 dido
X8 VDD VSS PCHG WREN SEL8 BL8 BL_8 DW8 DW_8 DR8 DR_8 dido
X9 VDD VSS PCHG WREN SEL9 BL9 BL_9 DW9 DW_9 DR9 DR_9 dido
X10 VDD VSS PCHG WREN SEL10 BL10 BL_10 DW10 DW_10 DR10 DR_10 dido
X11 VDD VSS PCHG WREN SEL11 BL11 BL_11 DW11 DW_11 DR11 DR_11 dido
X12 VDD VSS PCHG WREN SEL12 BL12 BL_12 DW12 DW_12 DR12 DR_12 dido
X13 VDD VSS PCHG WREN SEL13 BL13 BL_13 DW13 DW_13 DR13 DR_13 dido
X14 VDD VSS PCHG WREN SEL14 BL14 BL_14 DW14 DW_14 DR14 DR_14 dido
X15 VDD VSS PCHG WREN SEL15 BL15 BL_15 DW15 DW_15 DR15 DR_15 dido
X16 VDD VSS PCHG WREN SEL16 BL16 BL_16 DW16 DW_16 DR16 DR_16 dido
X17 VDD VSS PCHG WREN SEL17 BL17 BL_17 DW17 DW_17 DR17 DR_17 dido
X18 VDD VSS PCHG WREN SEL18 BL18 BL_18 DW18 DW_18 DR18 DR_18 dido
X19 VDD VSS PCHG WREN SEL19 BL19 BL_19 DW19 DW_19 DR19 DR_19 dido
X20 VDD VSS PCHG WREN SEL20 BL20 BL_20 DW20 DW_20 DR20 DR_20 dido
X21 VDD VSS PCHG WREN SEL21 BL21 BL_21 DW21 DW_21 DR21 DR_21 dido
X22 VDD VSS PCHG WREN SEL22 BL22 BL_22 DW22 DW_22 DR22 DR_22 dido
X23 VDD VSS PCHG WREN SEL23 BL23 BL_23 DW23 DW_23 DR23 DR_23 dido
X24 VDD VSS PCHG WREN SEL24 BL24 BL_24 DW24 DW_24 DR24 DR_24 dido
X25 VDD VSS PCHG WREN SEL25 BL25 BL_25 DW25 DW_25 DR25 DR_25 dido
X26 VDD VSS PCHG WREN SEL26 BL26 BL_26 DW26 DW_26 DR26 DR_26 dido
X27 VDD VSS PCHG WREN SEL27 BL27 BL_27 DW27 DW_27 DR27 DR_27 dido
X28 VDD VSS PCHG WREN SEL28 BL28 BL_28 DW28 DW_28 DR28 DR_28 dido
X29 VDD VSS PCHG WREN SEL29 BL29 BL_29 DW29 DW_29 DR29 DR_29 dido
X30 VDD VSS PCHG WREN SEL30 BL30 BL_30 DW30 DW_30 DR30 DR_30 dido
X31 VDD VSS PCHG WREN SEL31 BL31 BL_31 DW31 DW_31 DR31 DR_31 dido
X32 VDD VSS PCHG WREN SEL32 BL32 BL_32 DW32 DW_32 DR32 DR_32 dido
X33 VDD VSS PCHG WREN SEL33 BL33 BL_33 DW33 DW_33 DR33 DR_33 dido
X34 VDD VSS PCHG WREN SEL34 BL34 BL_34 DW34 DW_34 DR34 DR_34 dido
X35 VDD VSS PCHG WREN SEL35 BL35 BL_35 DW35 DW_35 DR35 DR_35 dido
X36 VDD VSS PCHG WREN SEL36 BL36 BL_36 DW36 DW_36 DR36 DR_36 dido
X37 VDD VSS PCHG WREN SEL37 BL37 BL_37 DW37 DW_37 DR37 DR_37 dido
X38 VDD VSS PCHG WREN SEL38 BL38 BL_38 DW38 DW_38 DR38 DR_38 dido
X39 VDD VSS PCHG WREN SEL39 BL39 BL_39 DW39 DW_39 DR39 DR_39 dido
X40 VDD VSS PCHG WREN SEL40 BL40 BL_40 DW40 DW_40 DR40 DR_40 dido
X41 VDD VSS PCHG WREN SEL41 BL41 BL_41 DW41 DW_41 DR41 DR_41 dido
X42 VDD VSS PCHG WREN SEL42 BL42 BL_42 DW42 DW_42 DR42 DR_42 dido
X43 VDD VSS PCHG WREN SEL43 BL43 BL_43 DW43 DW_43 DR43 DR_43 dido
X44 VDD VSS PCHG WREN SEL44 BL44 BL_44 DW44 DW_44 DR44 DR_44 dido
X45 VDD VSS PCHG WREN SEL45 BL45 BL_45 DW45 DW_45 DR45 DR_45 dido
X46 VDD VSS PCHG WREN SEL46 BL46 BL_46 DW46 DW_46 DR46 DR_46 dido
X47 VDD VSS PCHG WREN SEL47 BL47 BL_47 DW47 DW_47 DR47 DR_47 dido
X48 VDD VSS PCHG WREN SEL48 BL48 BL_48 DW48 DW_48 DR48 DR_48 dido
X49 VDD VSS PCHG WREN SEL49 BL49 BL_49 DW49 DW_49 DR49 DR_49 dido
X50 VDD VSS PCHG WREN SEL50 BL50 BL_50 DW50 DW_50 DR50 DR_50 dido
X51 VDD VSS PCHG WREN SEL51 BL51 BL_51 DW51 DW_51 DR51 DR_51 dido
X52 VDD VSS PCHG WREN SEL52 BL52 BL_52 DW52 DW_52 DR52 DR_52 dido
X53 VDD VSS PCHG WREN SEL53 BL53 BL_53 DW53 DW_53 DR53 DR_53 dido
X54 VDD VSS PCHG WREN SEL54 BL54 BL_54 DW54 DW_54 DR54 DR_54 dido
X55 VDD VSS PCHG WREN SEL55 BL55 BL_55 DW55 DW_55 DR55 DR_55 dido
X56 VDD VSS PCHG WREN SEL56 BL56 BL_56 DW56 DW_56 DR56 DR_56 dido
X57 VDD VSS PCHG WREN SEL57 BL57 BL_57 DW57 DW_57 DR57 DR_57 dido
X58 VDD VSS PCHG WREN SEL58 BL58 BL_58 DW58 DW_58 DR58 DR_58 dido
X59 VDD VSS PCHG WREN SEL59 BL59 BL_59 DW59 DW_59 DR59 DR_59 dido
X60 VDD VSS PCHG WREN SEL60 BL60 BL_60 DW60 DW_60 DR60 DR_60 dido
X61 VDD VSS PCHG WREN SEL61 BL61 BL_61 DW61 DW_61 DR61 DR_61 dido
X62 VDD VSS PCHG WREN SEL62 BL62 BL_62 DW62 DW_62 DR62 DR_62 dido
X63 VDD VSS PCHG WREN SEL63 BL63 BL_63 DW63 DW_63 DR63 DR_63 dido
X64 VDD VSS PCHG WREN SEL64 BL64 BL_64 DW64 DW_64 DR64 DR_64 dido
X65 VDD VSS PCHG WREN SEL65 BL65 BL_65 DW65 DW_65 DR65 DR_65 dido
X66 VDD VSS PCHG WREN SEL66 BL66 BL_66 DW66 DW_66 DR66 DR_66 dido
X67 VDD VSS PCHG WREN SEL67 BL67 BL_67 DW67 DW_67 DR67 DR_67 dido
X68 VDD VSS PCHG WREN SEL68 BL68 BL_68 DW68 DW_68 DR68 DR_68 dido
X69 VDD VSS PCHG WREN SEL69 BL69 BL_69 DW69 DW_69 DR69 DR_69 dido
X70 VDD VSS PCHG WREN SEL70 BL70 BL_70 DW70 DW_70 DR70 DR_70 dido
X71 VDD VSS PCHG WREN SEL71 BL71 BL_71 DW71 DW_71 DR71 DR_71 dido
X72 VDD VSS PCHG WREN SEL72 BL72 BL_72 DW72 DW_72 DR72 DR_72 dido
X73 VDD VSS PCHG WREN SEL73 BL73 BL_73 DW73 DW_73 DR73 DR_73 dido
X74 VDD VSS PCHG WREN SEL74 BL74 BL_74 DW74 DW_74 DR74 DR_74 dido
X75 VDD VSS PCHG WREN SEL75 BL75 BL_75 DW75 DW_75 DR75 DR_75 dido
X76 VDD VSS PCHG WREN SEL76 BL76 BL_76 DW76 DW_76 DR76 DR_76 dido
X77 VDD VSS PCHG WREN SEL77 BL77 BL_77 DW77 DW_77 DR77 DR_77 dido
X78 VDD VSS PCHG WREN SEL78 BL78 BL_78 DW78 DW_78 DR78 DR_78 dido
X79 VDD VSS PCHG WREN SEL79 BL79 BL_79 DW79 DW_79 DR79 DR_79 dido
X80 VDD VSS PCHG WREN SEL80 BL80 BL_80 DW80 DW_80 DR80 DR_80 dido
X81 VDD VSS PCHG WREN SEL81 BL81 BL_81 DW81 DW_81 DR81 DR_81 dido
X82 VDD VSS PCHG WREN SEL82 BL82 BL_82 DW82 DW_82 DR82 DR_82 dido
X83 VDD VSS PCHG WREN SEL83 BL83 BL_83 DW83 DW_83 DR83 DR_83 dido
X84 VDD VSS PCHG WREN SEL84 BL84 BL_84 DW84 DW_84 DR84 DR_84 dido
X85 VDD VSS PCHG WREN SEL85 BL85 BL_85 DW85 DW_85 DR85 DR_85 dido
X86 VDD VSS PCHG WREN SEL86 BL86 BL_86 DW86 DW_86 DR86 DR_86 dido
X87 VDD VSS PCHG WREN SEL87 BL87 BL_87 DW87 DW_87 DR87 DR_87 dido
X88 VDD VSS PCHG WREN SEL88 BL88 BL_88 DW88 DW_88 DR88 DR_88 dido
X89 VDD VSS PCHG WREN SEL89 BL89 BL_89 DW89 DW_89 DR89 DR_89 dido
X90 VDD VSS PCHG WREN SEL90 BL90 BL_90 DW90 DW_90 DR90 DR_90 dido
X91 VDD VSS PCHG WREN SEL91 BL91 BL_91 DW91 DW_91 DR91 DR_91 dido
X92 VDD VSS PCHG WREN SEL92 BL92 BL_92 DW92 DW_92 DR92 DR_92 dido
X93 VDD VSS PCHG WREN SEL93 BL93 BL_93 DW93 DW_93 DR93 DR_93 dido
X94 VDD VSS PCHG WREN SEL94 BL94 BL_94 DW94 DW_94 DR94 DR_94 dido
X95 VDD VSS PCHG WREN SEL95 BL95 BL_95 DW95 DW_95 DR95 DR_95 dido
X96 VDD VSS PCHG WREN SEL96 BL96 BL_96 DW96 DW_96 DR96 DR_96 dido
X97 VDD VSS PCHG WREN SEL97 BL97 BL_97 DW97 DW_97 DR97 DR_97 dido
X98 VDD VSS PCHG WREN SEL98 BL98 BL_98 DW98 DW_98 DR98 DR_98 dido
X99 VDD VSS PCHG WREN SEL99 BL99 BL_99 DW99 DW_99 DR99 DR_99 dido
X100 VDD VSS PCHG WREN SEL100 BL100 BL_100 DW100 DW_100 DR100 DR_100 dido
X101 VDD VSS PCHG WREN SEL101 BL101 BL_101 DW101 DW_101 DR101 DR_101 dido
X102 VDD VSS PCHG WREN SEL102 BL102 BL_102 DW102 DW_102 DR102 DR_102 dido
X103 VDD VSS PCHG WREN SEL103 BL103 BL_103 DW103 DW_103 DR103 DR_103 dido
X104 VDD VSS PCHG WREN SEL104 BL104 BL_104 DW104 DW_104 DR104 DR_104 dido
X105 VDD VSS PCHG WREN SEL105 BL105 BL_105 DW105 DW_105 DR105 DR_105 dido
X106 VDD VSS PCHG WREN SEL106 BL106 BL_106 DW106 DW_106 DR106 DR_106 dido
X107 VDD VSS PCHG WREN SEL107 BL107 BL_107 DW107 DW_107 DR107 DR_107 dido
X108 VDD VSS PCHG WREN SEL108 BL108 BL_108 DW108 DW_108 DR108 DR_108 dido
X109 VDD VSS PCHG WREN SEL109 BL109 BL_109 DW109 DW_109 DR109 DR_109 dido
X110 VDD VSS PCHG WREN SEL110 BL110 BL_110 DW110 DW_110 DR110 DR_110 dido
X111 VDD VSS PCHG WREN SEL111 BL111 BL_111 DW111 DW_111 DR111 DR_111 dido
X112 VDD VSS PCHG WREN SEL112 BL112 BL_112 DW112 DW_112 DR112 DR_112 dido
X113 VDD VSS PCHG WREN SEL113 BL113 BL_113 DW113 DW_113 DR113 DR_113 dido
X114 VDD VSS PCHG WREN SEL114 BL114 BL_114 DW114 DW_114 DR114 DR_114 dido
X115 VDD VSS PCHG WREN SEL115 BL115 BL_115 DW115 DW_115 DR115 DR_115 dido
X116 VDD VSS PCHG WREN SEL116 BL116 BL_116 DW116 DW_116 DR116 DR_116 dido
X117 VDD VSS PCHG WREN SEL117 BL117 BL_117 DW117 DW_117 DR117 DR_117 dido
X118 VDD VSS PCHG WREN SEL118 BL118 BL_118 DW118 DW_118 DR118 DR_118 dido
X119 VDD VSS PCHG WREN SEL119 BL119 BL_119 DW119 DW_119 DR119 DR_119 dido
X120 VDD VSS PCHG WREN SEL120 BL120 BL_120 DW120 DW_120 DR120 DR_120 dido
X121 VDD VSS PCHG WREN SEL121 BL121 BL_121 DW121 DW_121 DR121 DR_121 dido
X122 VDD VSS PCHG WREN SEL122 BL122 BL_122 DW122 DW_122 DR122 DR_122 dido
X123 VDD VSS PCHG WREN SEL123 BL123 BL_123 DW123 DW_123 DR123 DR_123 dido
X124 VDD VSS PCHG WREN SEL124 BL124 BL_124 DW124 DW_124 DR124 DR_124 dido
X125 VDD VSS PCHG WREN SEL125 BL125 BL_125 DW125 DW_125 DR125 DR_125 dido
X126 VDD VSS PCHG WREN SEL126 BL126 BL_126 DW126 DW_126 DR126 DR_126 dido
X127 VDD VSS PCHG WREN SEL127 BL127 BL_127 DW127 DW_127 DR127 DR_127 dido
X128 VDD VSS PCHG WREN SEL128 BL128 BL_128 DW128 DW_128 DR128 DR_128 dido
X129 VDD VSS PCHG WREN SEL129 BL129 BL_129 DW129 DW_129 DR129 DR_129 dido
X130 VDD VSS PCHG WREN SEL130 BL130 BL_130 DW130 DW_130 DR130 DR_130 dido
X131 VDD VSS PCHG WREN SEL131 BL131 BL_131 DW131 DW_131 DR131 DR_131 dido
X132 VDD VSS PCHG WREN SEL132 BL132 BL_132 DW132 DW_132 DR132 DR_132 dido
X133 VDD VSS PCHG WREN SEL133 BL133 BL_133 DW133 DW_133 DR133 DR_133 dido
X134 VDD VSS PCHG WREN SEL134 BL134 BL_134 DW134 DW_134 DR134 DR_134 dido
X135 VDD VSS PCHG WREN SEL135 BL135 BL_135 DW135 DW_135 DR135 DR_135 dido
X136 VDD VSS PCHG WREN SEL136 BL136 BL_136 DW136 DW_136 DR136 DR_136 dido
X137 VDD VSS PCHG WREN SEL137 BL137 BL_137 DW137 DW_137 DR137 DR_137 dido
X138 VDD VSS PCHG WREN SEL138 BL138 BL_138 DW138 DW_138 DR138 DR_138 dido
X139 VDD VSS PCHG WREN SEL139 BL139 BL_139 DW139 DW_139 DR139 DR_139 dido
X140 VDD VSS PCHG WREN SEL140 BL140 BL_140 DW140 DW_140 DR140 DR_140 dido
X141 VDD VSS PCHG WREN SEL141 BL141 BL_141 DW141 DW_141 DR141 DR_141 dido
X142 VDD VSS PCHG WREN SEL142 BL142 BL_142 DW142 DW_142 DR142 DR_142 dido
X143 VDD VSS PCHG WREN SEL143 BL143 BL_143 DW143 DW_143 DR143 DR_143 dido
X144 VDD VSS PCHG WREN SEL144 BL144 BL_144 DW144 DW_144 DR144 DR_144 dido
X145 VDD VSS PCHG WREN SEL145 BL145 BL_145 DW145 DW_145 DR145 DR_145 dido
X146 VDD VSS PCHG WREN SEL146 BL146 BL_146 DW146 DW_146 DR146 DR_146 dido
X147 VDD VSS PCHG WREN SEL147 BL147 BL_147 DW147 DW_147 DR147 DR_147 dido
X148 VDD VSS PCHG WREN SEL148 BL148 BL_148 DW148 DW_148 DR148 DR_148 dido
X149 VDD VSS PCHG WREN SEL149 BL149 BL_149 DW149 DW_149 DR149 DR_149 dido
X150 VDD VSS PCHG WREN SEL150 BL150 BL_150 DW150 DW_150 DR150 DR_150 dido
X151 VDD VSS PCHG WREN SEL151 BL151 BL_151 DW151 DW_151 DR151 DR_151 dido
X152 VDD VSS PCHG WREN SEL152 BL152 BL_152 DW152 DW_152 DR152 DR_152 dido
X153 VDD VSS PCHG WREN SEL153 BL153 BL_153 DW153 DW_153 DR153 DR_153 dido
X154 VDD VSS PCHG WREN SEL154 BL154 BL_154 DW154 DW_154 DR154 DR_154 dido
X155 VDD VSS PCHG WREN SEL155 BL155 BL_155 DW155 DW_155 DR155 DR_155 dido
X156 VDD VSS PCHG WREN SEL156 BL156 BL_156 DW156 DW_156 DR156 DR_156 dido
X157 VDD VSS PCHG WREN SEL157 BL157 BL_157 DW157 DW_157 DR157 DR_157 dido
X158 VDD VSS PCHG WREN SEL158 BL158 BL_158 DW158 DW_158 DR158 DR_158 dido
X159 VDD VSS PCHG WREN SEL159 BL159 BL_159 DW159 DW_159 DR159 DR_159 dido
X160 VDD VSS PCHG WREN SEL160 BL160 BL_160 DW160 DW_160 DR160 DR_160 dido
X161 VDD VSS PCHG WREN SEL161 BL161 BL_161 DW161 DW_161 DR161 DR_161 dido
X162 VDD VSS PCHG WREN SEL162 BL162 BL_162 DW162 DW_162 DR162 DR_162 dido
X163 VDD VSS PCHG WREN SEL163 BL163 BL_163 DW163 DW_163 DR163 DR_163 dido
X164 VDD VSS PCHG WREN SEL164 BL164 BL_164 DW164 DW_164 DR164 DR_164 dido
X165 VDD VSS PCHG WREN SEL165 BL165 BL_165 DW165 DW_165 DR165 DR_165 dido
X166 VDD VSS PCHG WREN SEL166 BL166 BL_166 DW166 DW_166 DR166 DR_166 dido
X167 VDD VSS PCHG WREN SEL167 BL167 BL_167 DW167 DW_167 DR167 DR_167 dido
X168 VDD VSS PCHG WREN SEL168 BL168 BL_168 DW168 DW_168 DR168 DR_168 dido
X169 VDD VSS PCHG WREN SEL169 BL169 BL_169 DW169 DW_169 DR169 DR_169 dido
X170 VDD VSS PCHG WREN SEL170 BL170 BL_170 DW170 DW_170 DR170 DR_170 dido
X171 VDD VSS PCHG WREN SEL171 BL171 BL_171 DW171 DW_171 DR171 DR_171 dido
X172 VDD VSS PCHG WREN SEL172 BL172 BL_172 DW172 DW_172 DR172 DR_172 dido
X173 VDD VSS PCHG WREN SEL173 BL173 BL_173 DW173 DW_173 DR173 DR_173 dido
X174 VDD VSS PCHG WREN SEL174 BL174 BL_174 DW174 DW_174 DR174 DR_174 dido
X175 VDD VSS PCHG WREN SEL175 BL175 BL_175 DW175 DW_175 DR175 DR_175 dido
X176 VDD VSS PCHG WREN SEL176 BL176 BL_176 DW176 DW_176 DR176 DR_176 dido
X177 VDD VSS PCHG WREN SEL177 BL177 BL_177 DW177 DW_177 DR177 DR_177 dido
X178 VDD VSS PCHG WREN SEL178 BL178 BL_178 DW178 DW_178 DR178 DR_178 dido
X179 VDD VSS PCHG WREN SEL179 BL179 BL_179 DW179 DW_179 DR179 DR_179 dido
X180 VDD VSS PCHG WREN SEL180 BL180 BL_180 DW180 DW_180 DR180 DR_180 dido
X181 VDD VSS PCHG WREN SEL181 BL181 BL_181 DW181 DW_181 DR181 DR_181 dido
X182 VDD VSS PCHG WREN SEL182 BL182 BL_182 DW182 DW_182 DR182 DR_182 dido
X183 VDD VSS PCHG WREN SEL183 BL183 BL_183 DW183 DW_183 DR183 DR_183 dido
X184 VDD VSS PCHG WREN SEL184 BL184 BL_184 DW184 DW_184 DR184 DR_184 dido
X185 VDD VSS PCHG WREN SEL185 BL185 BL_185 DW185 DW_185 DR185 DR_185 dido
X186 VDD VSS PCHG WREN SEL186 BL186 BL_186 DW186 DW_186 DR186 DR_186 dido
X187 VDD VSS PCHG WREN SEL187 BL187 BL_187 DW187 DW_187 DR187 DR_187 dido
X188 VDD VSS PCHG WREN SEL188 BL188 BL_188 DW188 DW_188 DR188 DR_188 dido
X189 VDD VSS PCHG WREN SEL189 BL189 BL_189 DW189 DW_189 DR189 DR_189 dido
X190 VDD VSS PCHG WREN SEL190 BL190 BL_190 DW190 DW_190 DR190 DR_190 dido
X191 VDD VSS PCHG WREN SEL191 BL191 BL_191 DW191 DW_191 DR191 DR_191 dido
X192 VDD VSS PCHG WREN SEL192 BL192 BL_192 DW192 DW_192 DR192 DR_192 dido
X193 VDD VSS PCHG WREN SEL193 BL193 BL_193 DW193 DW_193 DR193 DR_193 dido
X194 VDD VSS PCHG WREN SEL194 BL194 BL_194 DW194 DW_194 DR194 DR_194 dido
X195 VDD VSS PCHG WREN SEL195 BL195 BL_195 DW195 DW_195 DR195 DR_195 dido
X196 VDD VSS PCHG WREN SEL196 BL196 BL_196 DW196 DW_196 DR196 DR_196 dido
X197 VDD VSS PCHG WREN SEL197 BL197 BL_197 DW197 DW_197 DR197 DR_197 dido
X198 VDD VSS PCHG WREN SEL198 BL198 BL_198 DW198 DW_198 DR198 DR_198 dido
X199 VDD VSS PCHG WREN SEL199 BL199 BL_199 DW199 DW_199 DR199 DR_199 dido
X200 VDD VSS PCHG WREN SEL200 BL200 BL_200 DW200 DW_200 DR200 DR_200 dido
X201 VDD VSS PCHG WREN SEL201 BL201 BL_201 DW201 DW_201 DR201 DR_201 dido
X202 VDD VSS PCHG WREN SEL202 BL202 BL_202 DW202 DW_202 DR202 DR_202 dido
X203 VDD VSS PCHG WREN SEL203 BL203 BL_203 DW203 DW_203 DR203 DR_203 dido
X204 VDD VSS PCHG WREN SEL204 BL204 BL_204 DW204 DW_204 DR204 DR_204 dido
X205 VDD VSS PCHG WREN SEL205 BL205 BL_205 DW205 DW_205 DR205 DR_205 dido
X206 VDD VSS PCHG WREN SEL206 BL206 BL_206 DW206 DW_206 DR206 DR_206 dido
X207 VDD VSS PCHG WREN SEL207 BL207 BL_207 DW207 DW_207 DR207 DR_207 dido
X208 VDD VSS PCHG WREN SEL208 BL208 BL_208 DW208 DW_208 DR208 DR_208 dido
X209 VDD VSS PCHG WREN SEL209 BL209 BL_209 DW209 DW_209 DR209 DR_209 dido
X210 VDD VSS PCHG WREN SEL210 BL210 BL_210 DW210 DW_210 DR210 DR_210 dido
X211 VDD VSS PCHG WREN SEL211 BL211 BL_211 DW211 DW_211 DR211 DR_211 dido
X212 VDD VSS PCHG WREN SEL212 BL212 BL_212 DW212 DW_212 DR212 DR_212 dido
X213 VDD VSS PCHG WREN SEL213 BL213 BL_213 DW213 DW_213 DR213 DR_213 dido
X214 VDD VSS PCHG WREN SEL214 BL214 BL_214 DW214 DW_214 DR214 DR_214 dido
X215 VDD VSS PCHG WREN SEL215 BL215 BL_215 DW215 DW_215 DR215 DR_215 dido
X216 VDD VSS PCHG WREN SEL216 BL216 BL_216 DW216 DW_216 DR216 DR_216 dido
X217 VDD VSS PCHG WREN SEL217 BL217 BL_217 DW217 DW_217 DR217 DR_217 dido
X218 VDD VSS PCHG WREN SEL218 BL218 BL_218 DW218 DW_218 DR218 DR_218 dido
X219 VDD VSS PCHG WREN SEL219 BL219 BL_219 DW219 DW_219 DR219 DR_219 dido
X220 VDD VSS PCHG WREN SEL220 BL220 BL_220 DW220 DW_220 DR220 DR_220 dido
X221 VDD VSS PCHG WREN SEL221 BL221 BL_221 DW221 DW_221 DR221 DR_221 dido
X222 VDD VSS PCHG WREN SEL222 BL222 BL_222 DW222 DW_222 DR222 DR_222 dido
X223 VDD VSS PCHG WREN SEL223 BL223 BL_223 DW223 DW_223 DR223 DR_223 dido
X224 VDD VSS PCHG WREN SEL224 BL224 BL_224 DW224 DW_224 DR224 DR_224 dido
X225 VDD VSS PCHG WREN SEL225 BL225 BL_225 DW225 DW_225 DR225 DR_225 dido
X226 VDD VSS PCHG WREN SEL226 BL226 BL_226 DW226 DW_226 DR226 DR_226 dido
X227 VDD VSS PCHG WREN SEL227 BL227 BL_227 DW227 DW_227 DR227 DR_227 dido
X228 VDD VSS PCHG WREN SEL228 BL228 BL_228 DW228 DW_228 DR228 DR_228 dido
X229 VDD VSS PCHG WREN SEL229 BL229 BL_229 DW229 DW_229 DR229 DR_229 dido
X230 VDD VSS PCHG WREN SEL230 BL230 BL_230 DW230 DW_230 DR230 DR_230 dido
X231 VDD VSS PCHG WREN SEL231 BL231 BL_231 DW231 DW_231 DR231 DR_231 dido
X232 VDD VSS PCHG WREN SEL232 BL232 BL_232 DW232 DW_232 DR232 DR_232 dido
X233 VDD VSS PCHG WREN SEL233 BL233 BL_233 DW233 DW_233 DR233 DR_233 dido
X234 VDD VSS PCHG WREN SEL234 BL234 BL_234 DW234 DW_234 DR234 DR_234 dido
X235 VDD VSS PCHG WREN SEL235 BL235 BL_235 DW235 DW_235 DR235 DR_235 dido
X236 VDD VSS PCHG WREN SEL236 BL236 BL_236 DW236 DW_236 DR236 DR_236 dido
X237 VDD VSS PCHG WREN SEL237 BL237 BL_237 DW237 DW_237 DR237 DR_237 dido
X238 VDD VSS PCHG WREN SEL238 BL238 BL_238 DW238 DW_238 DR238 DR_238 dido
X239 VDD VSS PCHG WREN SEL239 BL239 BL_239 DW239 DW_239 DR239 DR_239 dido
X240 VDD VSS PCHG WREN SEL240 BL240 BL_240 DW240 DW_240 DR240 DR_240 dido
X241 VDD VSS PCHG WREN SEL241 BL241 BL_241 DW241 DW_241 DR241 DR_241 dido
X242 VDD VSS PCHG WREN SEL242 BL242 BL_242 DW242 DW_242 DR242 DR_242 dido
X243 VDD VSS PCHG WREN SEL243 BL243 BL_243 DW243 DW_243 DR243 DR_243 dido
X244 VDD VSS PCHG WREN SEL244 BL244 BL_244 DW244 DW_244 DR244 DR_244 dido
X245 VDD VSS PCHG WREN SEL245 BL245 BL_245 DW245 DW_245 DR245 DR_245 dido
X246 VDD VSS PCHG WREN SEL246 BL246 BL_246 DW246 DW_246 DR246 DR_246 dido
X247 VDD VSS PCHG WREN SEL247 BL247 BL_247 DW247 DW_247 DR247 DR_247 dido
X248 VDD VSS PCHG WREN SEL248 BL248 BL_248 DW248 DW_248 DR248 DR_248 dido
X249 VDD VSS PCHG WREN SEL249 BL249 BL_249 DW249 DW_249 DR249 DR_249 dido
X250 VDD VSS PCHG WREN SEL250 BL250 BL_250 DW250 DW_250 DR250 DR_250 dido
X251 VDD VSS PCHG WREN SEL251 BL251 BL_251 DW251 DW_251 DR251 DR_251 dido
X252 VDD VSS PCHG WREN SEL252 BL252 BL_252 DW252 DW_252 DR252 DR_252 dido
X253 VDD VSS PCHG WREN SEL253 BL253 BL_253 DW253 DW_253 DR253 DR_253 dido
X254 VDD VSS PCHG WREN SEL254 BL254 BL_254 DW254 DW_254 DR254 DR_254 dido
X255 VDD VSS PCHG WREN SEL255 BL255 BL_255 DW255 DW_255 DR255 DR_255 dido
X256 VDD VSS PCHG WREN SEL256 BL256 BL_256 DW256 DW_256 DR256 DR_256 dido
X257 VDD VSS PCHG WREN SEL257 BL257 BL_257 DW257 DW_257 DR257 DR_257 dido
X258 VDD VSS PCHG WREN SEL258 BL258 BL_258 DW258 DW_258 DR258 DR_258 dido
X259 VDD VSS PCHG WREN SEL259 BL259 BL_259 DW259 DW_259 DR259 DR_259 dido
X260 VDD VSS PCHG WREN SEL260 BL260 BL_260 DW260 DW_260 DR260 DR_260 dido
X261 VDD VSS PCHG WREN SEL261 BL261 BL_261 DW261 DW_261 DR261 DR_261 dido
X262 VDD VSS PCHG WREN SEL262 BL262 BL_262 DW262 DW_262 DR262 DR_262 dido
X263 VDD VSS PCHG WREN SEL263 BL263 BL_263 DW263 DW_263 DR263 DR_263 dido
X264 VDD VSS PCHG WREN SEL264 BL264 BL_264 DW264 DW_264 DR264 DR_264 dido
X265 VDD VSS PCHG WREN SEL265 BL265 BL_265 DW265 DW_265 DR265 DR_265 dido
X266 VDD VSS PCHG WREN SEL266 BL266 BL_266 DW266 DW_266 DR266 DR_266 dido
X267 VDD VSS PCHG WREN SEL267 BL267 BL_267 DW267 DW_267 DR267 DR_267 dido
X268 VDD VSS PCHG WREN SEL268 BL268 BL_268 DW268 DW_268 DR268 DR_268 dido
X269 VDD VSS PCHG WREN SEL269 BL269 BL_269 DW269 DW_269 DR269 DR_269 dido
X270 VDD VSS PCHG WREN SEL270 BL270 BL_270 DW270 DW_270 DR270 DR_270 dido
X271 VDD VSS PCHG WREN SEL271 BL271 BL_271 DW271 DW_271 DR271 DR_271 dido
X272 VDD VSS PCHG WREN SEL272 BL272 BL_272 DW272 DW_272 DR272 DR_272 dido
X273 VDD VSS PCHG WREN SEL273 BL273 BL_273 DW273 DW_273 DR273 DR_273 dido
X274 VDD VSS PCHG WREN SEL274 BL274 BL_274 DW274 DW_274 DR274 DR_274 dido
X275 VDD VSS PCHG WREN SEL275 BL275 BL_275 DW275 DW_275 DR275 DR_275 dido
X276 VDD VSS PCHG WREN SEL276 BL276 BL_276 DW276 DW_276 DR276 DR_276 dido
X277 VDD VSS PCHG WREN SEL277 BL277 BL_277 DW277 DW_277 DR277 DR_277 dido
X278 VDD VSS PCHG WREN SEL278 BL278 BL_278 DW278 DW_278 DR278 DR_278 dido
X279 VDD VSS PCHG WREN SEL279 BL279 BL_279 DW279 DW_279 DR279 DR_279 dido
X280 VDD VSS PCHG WREN SEL280 BL280 BL_280 DW280 DW_280 DR280 DR_280 dido
X281 VDD VSS PCHG WREN SEL281 BL281 BL_281 DW281 DW_281 DR281 DR_281 dido
X282 VDD VSS PCHG WREN SEL282 BL282 BL_282 DW282 DW_282 DR282 DR_282 dido
X283 VDD VSS PCHG WREN SEL283 BL283 BL_283 DW283 DW_283 DR283 DR_283 dido
X284 VDD VSS PCHG WREN SEL284 BL284 BL_284 DW284 DW_284 DR284 DR_284 dido
X285 VDD VSS PCHG WREN SEL285 BL285 BL_285 DW285 DW_285 DR285 DR_285 dido
X286 VDD VSS PCHG WREN SEL286 BL286 BL_286 DW286 DW_286 DR286 DR_286 dido
X287 VDD VSS PCHG WREN SEL287 BL287 BL_287 DW287 DW_287 DR287 DR_287 dido
X288 VDD VSS PCHG WREN SEL288 BL288 BL_288 DW288 DW_288 DR288 DR_288 dido
X289 VDD VSS PCHG WREN SEL289 BL289 BL_289 DW289 DW_289 DR289 DR_289 dido
X290 VDD VSS PCHG WREN SEL290 BL290 BL_290 DW290 DW_290 DR290 DR_290 dido
X291 VDD VSS PCHG WREN SEL291 BL291 BL_291 DW291 DW_291 DR291 DR_291 dido
X292 VDD VSS PCHG WREN SEL292 BL292 BL_292 DW292 DW_292 DR292 DR_292 dido
X293 VDD VSS PCHG WREN SEL293 BL293 BL_293 DW293 DW_293 DR293 DR_293 dido
X294 VDD VSS PCHG WREN SEL294 BL294 BL_294 DW294 DW_294 DR294 DR_294 dido
X295 VDD VSS PCHG WREN SEL295 BL295 BL_295 DW295 DW_295 DR295 DR_295 dido
X296 VDD VSS PCHG WREN SEL296 BL296 BL_296 DW296 DW_296 DR296 DR_296 dido
X297 VDD VSS PCHG WREN SEL297 BL297 BL_297 DW297 DW_297 DR297 DR_297 dido
X298 VDD VSS PCHG WREN SEL298 BL298 BL_298 DW298 DW_298 DR298 DR_298 dido
X299 VDD VSS PCHG WREN SEL299 BL299 BL_299 DW299 DW_299 DR299 DR_299 dido
X300 VDD VSS PCHG WREN SEL300 BL300 BL_300 DW300 DW_300 DR300 DR_300 dido
X301 VDD VSS PCHG WREN SEL301 BL301 BL_301 DW301 DW_301 DR301 DR_301 dido
X302 VDD VSS PCHG WREN SEL302 BL302 BL_302 DW302 DW_302 DR302 DR_302 dido
X303 VDD VSS PCHG WREN SEL303 BL303 BL_303 DW303 DW_303 DR303 DR_303 dido
X304 VDD VSS PCHG WREN SEL304 BL304 BL_304 DW304 DW_304 DR304 DR_304 dido
X305 VDD VSS PCHG WREN SEL305 BL305 BL_305 DW305 DW_305 DR305 DR_305 dido
X306 VDD VSS PCHG WREN SEL306 BL306 BL_306 DW306 DW_306 DR306 DR_306 dido
X307 VDD VSS PCHG WREN SEL307 BL307 BL_307 DW307 DW_307 DR307 DR_307 dido
X308 VDD VSS PCHG WREN SEL308 BL308 BL_308 DW308 DW_308 DR308 DR_308 dido
X309 VDD VSS PCHG WREN SEL309 BL309 BL_309 DW309 DW_309 DR309 DR_309 dido
X310 VDD VSS PCHG WREN SEL310 BL310 BL_310 DW310 DW_310 DR310 DR_310 dido
X311 VDD VSS PCHG WREN SEL311 BL311 BL_311 DW311 DW_311 DR311 DR_311 dido
X312 VDD VSS PCHG WREN SEL312 BL312 BL_312 DW312 DW_312 DR312 DR_312 dido
X313 VDD VSS PCHG WREN SEL313 BL313 BL_313 DW313 DW_313 DR313 DR_313 dido
X314 VDD VSS PCHG WREN SEL314 BL314 BL_314 DW314 DW_314 DR314 DR_314 dido
X315 VDD VSS PCHG WREN SEL315 BL315 BL_315 DW315 DW_315 DR315 DR_315 dido
X316 VDD VSS PCHG WREN SEL316 BL316 BL_316 DW316 DW_316 DR316 DR_316 dido
X317 VDD VSS PCHG WREN SEL317 BL317 BL_317 DW317 DW_317 DR317 DR_317 dido
X318 VDD VSS PCHG WREN SEL318 BL318 BL_318 DW318 DW_318 DR318 DR_318 dido
X319 VDD VSS PCHG WREN SEL319 BL319 BL_319 DW319 DW_319 DR319 DR_319 dido
X320 VDD VSS PCHG WREN SEL320 BL320 BL_320 DW320 DW_320 DR320 DR_320 dido
X321 VDD VSS PCHG WREN SEL321 BL321 BL_321 DW321 DW_321 DR321 DR_321 dido
X322 VDD VSS PCHG WREN SEL322 BL322 BL_322 DW322 DW_322 DR322 DR_322 dido
X323 VDD VSS PCHG WREN SEL323 BL323 BL_323 DW323 DW_323 DR323 DR_323 dido
X324 VDD VSS PCHG WREN SEL324 BL324 BL_324 DW324 DW_324 DR324 DR_324 dido
X325 VDD VSS PCHG WREN SEL325 BL325 BL_325 DW325 DW_325 DR325 DR_325 dido
X326 VDD VSS PCHG WREN SEL326 BL326 BL_326 DW326 DW_326 DR326 DR_326 dido
X327 VDD VSS PCHG WREN SEL327 BL327 BL_327 DW327 DW_327 DR327 DR_327 dido
X328 VDD VSS PCHG WREN SEL328 BL328 BL_328 DW328 DW_328 DR328 DR_328 dido
X329 VDD VSS PCHG WREN SEL329 BL329 BL_329 DW329 DW_329 DR329 DR_329 dido
X330 VDD VSS PCHG WREN SEL330 BL330 BL_330 DW330 DW_330 DR330 DR_330 dido
X331 VDD VSS PCHG WREN SEL331 BL331 BL_331 DW331 DW_331 DR331 DR_331 dido
X332 VDD VSS PCHG WREN SEL332 BL332 BL_332 DW332 DW_332 DR332 DR_332 dido
X333 VDD VSS PCHG WREN SEL333 BL333 BL_333 DW333 DW_333 DR333 DR_333 dido
X334 VDD VSS PCHG WREN SEL334 BL334 BL_334 DW334 DW_334 DR334 DR_334 dido
X335 VDD VSS PCHG WREN SEL335 BL335 BL_335 DW335 DW_335 DR335 DR_335 dido
X336 VDD VSS PCHG WREN SEL336 BL336 BL_336 DW336 DW_336 DR336 DR_336 dido
X337 VDD VSS PCHG WREN SEL337 BL337 BL_337 DW337 DW_337 DR337 DR_337 dido
X338 VDD VSS PCHG WREN SEL338 BL338 BL_338 DW338 DW_338 DR338 DR_338 dido
X339 VDD VSS PCHG WREN SEL339 BL339 BL_339 DW339 DW_339 DR339 DR_339 dido
X340 VDD VSS PCHG WREN SEL340 BL340 BL_340 DW340 DW_340 DR340 DR_340 dido
X341 VDD VSS PCHG WREN SEL341 BL341 BL_341 DW341 DW_341 DR341 DR_341 dido
X342 VDD VSS PCHG WREN SEL342 BL342 BL_342 DW342 DW_342 DR342 DR_342 dido
X343 VDD VSS PCHG WREN SEL343 BL343 BL_343 DW343 DW_343 DR343 DR_343 dido
X344 VDD VSS PCHG WREN SEL344 BL344 BL_344 DW344 DW_344 DR344 DR_344 dido
X345 VDD VSS PCHG WREN SEL345 BL345 BL_345 DW345 DW_345 DR345 DR_345 dido
X346 VDD VSS PCHG WREN SEL346 BL346 BL_346 DW346 DW_346 DR346 DR_346 dido
X347 VDD VSS PCHG WREN SEL347 BL347 BL_347 DW347 DW_347 DR347 DR_347 dido
X348 VDD VSS PCHG WREN SEL348 BL348 BL_348 DW348 DW_348 DR348 DR_348 dido
X349 VDD VSS PCHG WREN SEL349 BL349 BL_349 DW349 DW_349 DR349 DR_349 dido
X350 VDD VSS PCHG WREN SEL350 BL350 BL_350 DW350 DW_350 DR350 DR_350 dido
X351 VDD VSS PCHG WREN SEL351 BL351 BL_351 DW351 DW_351 DR351 DR_351 dido
X352 VDD VSS PCHG WREN SEL352 BL352 BL_352 DW352 DW_352 DR352 DR_352 dido
X353 VDD VSS PCHG WREN SEL353 BL353 BL_353 DW353 DW_353 DR353 DR_353 dido
X354 VDD VSS PCHG WREN SEL354 BL354 BL_354 DW354 DW_354 DR354 DR_354 dido
X355 VDD VSS PCHG WREN SEL355 BL355 BL_355 DW355 DW_355 DR355 DR_355 dido
X356 VDD VSS PCHG WREN SEL356 BL356 BL_356 DW356 DW_356 DR356 DR_356 dido
X357 VDD VSS PCHG WREN SEL357 BL357 BL_357 DW357 DW_357 DR357 DR_357 dido
X358 VDD VSS PCHG WREN SEL358 BL358 BL_358 DW358 DW_358 DR358 DR_358 dido
X359 VDD VSS PCHG WREN SEL359 BL359 BL_359 DW359 DW_359 DR359 DR_359 dido
X360 VDD VSS PCHG WREN SEL360 BL360 BL_360 DW360 DW_360 DR360 DR_360 dido
X361 VDD VSS PCHG WREN SEL361 BL361 BL_361 DW361 DW_361 DR361 DR_361 dido
X362 VDD VSS PCHG WREN SEL362 BL362 BL_362 DW362 DW_362 DR362 DR_362 dido
X363 VDD VSS PCHG WREN SEL363 BL363 BL_363 DW363 DW_363 DR363 DR_363 dido
X364 VDD VSS PCHG WREN SEL364 BL364 BL_364 DW364 DW_364 DR364 DR_364 dido
X365 VDD VSS PCHG WREN SEL365 BL365 BL_365 DW365 DW_365 DR365 DR_365 dido
X366 VDD VSS PCHG WREN SEL366 BL366 BL_366 DW366 DW_366 DR366 DR_366 dido
X367 VDD VSS PCHG WREN SEL367 BL367 BL_367 DW367 DW_367 DR367 DR_367 dido
X368 VDD VSS PCHG WREN SEL368 BL368 BL_368 DW368 DW_368 DR368 DR_368 dido
X369 VDD VSS PCHG WREN SEL369 BL369 BL_369 DW369 DW_369 DR369 DR_369 dido
X370 VDD VSS PCHG WREN SEL370 BL370 BL_370 DW370 DW_370 DR370 DR_370 dido
X371 VDD VSS PCHG WREN SEL371 BL371 BL_371 DW371 DW_371 DR371 DR_371 dido
X372 VDD VSS PCHG WREN SEL372 BL372 BL_372 DW372 DW_372 DR372 DR_372 dido
X373 VDD VSS PCHG WREN SEL373 BL373 BL_373 DW373 DW_373 DR373 DR_373 dido
X374 VDD VSS PCHG WREN SEL374 BL374 BL_374 DW374 DW_374 DR374 DR_374 dido
X375 VDD VSS PCHG WREN SEL375 BL375 BL_375 DW375 DW_375 DR375 DR_375 dido
X376 VDD VSS PCHG WREN SEL376 BL376 BL_376 DW376 DW_376 DR376 DR_376 dido
X377 VDD VSS PCHG WREN SEL377 BL377 BL_377 DW377 DW_377 DR377 DR_377 dido
X378 VDD VSS PCHG WREN SEL378 BL378 BL_378 DW378 DW_378 DR378 DR_378 dido
X379 VDD VSS PCHG WREN SEL379 BL379 BL_379 DW379 DW_379 DR379 DR_379 dido
X380 VDD VSS PCHG WREN SEL380 BL380 BL_380 DW380 DW_380 DR380 DR_380 dido
X381 VDD VSS PCHG WREN SEL381 BL381 BL_381 DW381 DW_381 DR381 DR_381 dido
X382 VDD VSS PCHG WREN SEL382 BL382 BL_382 DW382 DW_382 DR382 DR_382 dido
X383 VDD VSS PCHG WREN SEL383 BL383 BL_383 DW383 DW_383 DR383 DR_383 dido
X384 VDD VSS PCHG WREN SEL384 BL384 BL_384 DW384 DW_384 DR384 DR_384 dido
X385 VDD VSS PCHG WREN SEL385 BL385 BL_385 DW385 DW_385 DR385 DR_385 dido
X386 VDD VSS PCHG WREN SEL386 BL386 BL_386 DW386 DW_386 DR386 DR_386 dido
X387 VDD VSS PCHG WREN SEL387 BL387 BL_387 DW387 DW_387 DR387 DR_387 dido
X388 VDD VSS PCHG WREN SEL388 BL388 BL_388 DW388 DW_388 DR388 DR_388 dido
X389 VDD VSS PCHG WREN SEL389 BL389 BL_389 DW389 DW_389 DR389 DR_389 dido
X390 VDD VSS PCHG WREN SEL390 BL390 BL_390 DW390 DW_390 DR390 DR_390 dido
X391 VDD VSS PCHG WREN SEL391 BL391 BL_391 DW391 DW_391 DR391 DR_391 dido
X392 VDD VSS PCHG WREN SEL392 BL392 BL_392 DW392 DW_392 DR392 DR_392 dido
X393 VDD VSS PCHG WREN SEL393 BL393 BL_393 DW393 DW_393 DR393 DR_393 dido
X394 VDD VSS PCHG WREN SEL394 BL394 BL_394 DW394 DW_394 DR394 DR_394 dido
X395 VDD VSS PCHG WREN SEL395 BL395 BL_395 DW395 DW_395 DR395 DR_395 dido
X396 VDD VSS PCHG WREN SEL396 BL396 BL_396 DW396 DW_396 DR396 DR_396 dido
X397 VDD VSS PCHG WREN SEL397 BL397 BL_397 DW397 DW_397 DR397 DR_397 dido
X398 VDD VSS PCHG WREN SEL398 BL398 BL_398 DW398 DW_398 DR398 DR_398 dido
X399 VDD VSS PCHG WREN SEL399 BL399 BL_399 DW399 DW_399 DR399 DR_399 dido
X400 VDD VSS PCHG WREN SEL400 BL400 BL_400 DW400 DW_400 DR400 DR_400 dido
X401 VDD VSS PCHG WREN SEL401 BL401 BL_401 DW401 DW_401 DR401 DR_401 dido
X402 VDD VSS PCHG WREN SEL402 BL402 BL_402 DW402 DW_402 DR402 DR_402 dido
X403 VDD VSS PCHG WREN SEL403 BL403 BL_403 DW403 DW_403 DR403 DR_403 dido
X404 VDD VSS PCHG WREN SEL404 BL404 BL_404 DW404 DW_404 DR404 DR_404 dido
X405 VDD VSS PCHG WREN SEL405 BL405 BL_405 DW405 DW_405 DR405 DR_405 dido
X406 VDD VSS PCHG WREN SEL406 BL406 BL_406 DW406 DW_406 DR406 DR_406 dido
X407 VDD VSS PCHG WREN SEL407 BL407 BL_407 DW407 DW_407 DR407 DR_407 dido
X408 VDD VSS PCHG WREN SEL408 BL408 BL_408 DW408 DW_408 DR408 DR_408 dido
X409 VDD VSS PCHG WREN SEL409 BL409 BL_409 DW409 DW_409 DR409 DR_409 dido
X410 VDD VSS PCHG WREN SEL410 BL410 BL_410 DW410 DW_410 DR410 DR_410 dido
X411 VDD VSS PCHG WREN SEL411 BL411 BL_411 DW411 DW_411 DR411 DR_411 dido
X412 VDD VSS PCHG WREN SEL412 BL412 BL_412 DW412 DW_412 DR412 DR_412 dido
X413 VDD VSS PCHG WREN SEL413 BL413 BL_413 DW413 DW_413 DR413 DR_413 dido
X414 VDD VSS PCHG WREN SEL414 BL414 BL_414 DW414 DW_414 DR414 DR_414 dido
X415 VDD VSS PCHG WREN SEL415 BL415 BL_415 DW415 DW_415 DR415 DR_415 dido
X416 VDD VSS PCHG WREN SEL416 BL416 BL_416 DW416 DW_416 DR416 DR_416 dido
X417 VDD VSS PCHG WREN SEL417 BL417 BL_417 DW417 DW_417 DR417 DR_417 dido
X418 VDD VSS PCHG WREN SEL418 BL418 BL_418 DW418 DW_418 DR418 DR_418 dido
X419 VDD VSS PCHG WREN SEL419 BL419 BL_419 DW419 DW_419 DR419 DR_419 dido
X420 VDD VSS PCHG WREN SEL420 BL420 BL_420 DW420 DW_420 DR420 DR_420 dido
X421 VDD VSS PCHG WREN SEL421 BL421 BL_421 DW421 DW_421 DR421 DR_421 dido
X422 VDD VSS PCHG WREN SEL422 BL422 BL_422 DW422 DW_422 DR422 DR_422 dido
X423 VDD VSS PCHG WREN SEL423 BL423 BL_423 DW423 DW_423 DR423 DR_423 dido
X424 VDD VSS PCHG WREN SEL424 BL424 BL_424 DW424 DW_424 DR424 DR_424 dido
X425 VDD VSS PCHG WREN SEL425 BL425 BL_425 DW425 DW_425 DR425 DR_425 dido
X426 VDD VSS PCHG WREN SEL426 BL426 BL_426 DW426 DW_426 DR426 DR_426 dido
X427 VDD VSS PCHG WREN SEL427 BL427 BL_427 DW427 DW_427 DR427 DR_427 dido
X428 VDD VSS PCHG WREN SEL428 BL428 BL_428 DW428 DW_428 DR428 DR_428 dido
X429 VDD VSS PCHG WREN SEL429 BL429 BL_429 DW429 DW_429 DR429 DR_429 dido
X430 VDD VSS PCHG WREN SEL430 BL430 BL_430 DW430 DW_430 DR430 DR_430 dido
X431 VDD VSS PCHG WREN SEL431 BL431 BL_431 DW431 DW_431 DR431 DR_431 dido
X432 VDD VSS PCHG WREN SEL432 BL432 BL_432 DW432 DW_432 DR432 DR_432 dido
X433 VDD VSS PCHG WREN SEL433 BL433 BL_433 DW433 DW_433 DR433 DR_433 dido
X434 VDD VSS PCHG WREN SEL434 BL434 BL_434 DW434 DW_434 DR434 DR_434 dido
X435 VDD VSS PCHG WREN SEL435 BL435 BL_435 DW435 DW_435 DR435 DR_435 dido
X436 VDD VSS PCHG WREN SEL436 BL436 BL_436 DW436 DW_436 DR436 DR_436 dido
X437 VDD VSS PCHG WREN SEL437 BL437 BL_437 DW437 DW_437 DR437 DR_437 dido
X438 VDD VSS PCHG WREN SEL438 BL438 BL_438 DW438 DW_438 DR438 DR_438 dido
X439 VDD VSS PCHG WREN SEL439 BL439 BL_439 DW439 DW_439 DR439 DR_439 dido
X440 VDD VSS PCHG WREN SEL440 BL440 BL_440 DW440 DW_440 DR440 DR_440 dido
X441 VDD VSS PCHG WREN SEL441 BL441 BL_441 DW441 DW_441 DR441 DR_441 dido
X442 VDD VSS PCHG WREN SEL442 BL442 BL_442 DW442 DW_442 DR442 DR_442 dido
X443 VDD VSS PCHG WREN SEL443 BL443 BL_443 DW443 DW_443 DR443 DR_443 dido
X444 VDD VSS PCHG WREN SEL444 BL444 BL_444 DW444 DW_444 DR444 DR_444 dido
X445 VDD VSS PCHG WREN SEL445 BL445 BL_445 DW445 DW_445 DR445 DR_445 dido
X446 VDD VSS PCHG WREN SEL446 BL446 BL_446 DW446 DW_446 DR446 DR_446 dido
X447 VDD VSS PCHG WREN SEL447 BL447 BL_447 DW447 DW_447 DR447 DR_447 dido
X448 VDD VSS PCHG WREN SEL448 BL448 BL_448 DW448 DW_448 DR448 DR_448 dido
X449 VDD VSS PCHG WREN SEL449 BL449 BL_449 DW449 DW_449 DR449 DR_449 dido
X450 VDD VSS PCHG WREN SEL450 BL450 BL_450 DW450 DW_450 DR450 DR_450 dido
X451 VDD VSS PCHG WREN SEL451 BL451 BL_451 DW451 DW_451 DR451 DR_451 dido
X452 VDD VSS PCHG WREN SEL452 BL452 BL_452 DW452 DW_452 DR452 DR_452 dido
X453 VDD VSS PCHG WREN SEL453 BL453 BL_453 DW453 DW_453 DR453 DR_453 dido
X454 VDD VSS PCHG WREN SEL454 BL454 BL_454 DW454 DW_454 DR454 DR_454 dido
X455 VDD VSS PCHG WREN SEL455 BL455 BL_455 DW455 DW_455 DR455 DR_455 dido
X456 VDD VSS PCHG WREN SEL456 BL456 BL_456 DW456 DW_456 DR456 DR_456 dido
X457 VDD VSS PCHG WREN SEL457 BL457 BL_457 DW457 DW_457 DR457 DR_457 dido
X458 VDD VSS PCHG WREN SEL458 BL458 BL_458 DW458 DW_458 DR458 DR_458 dido
X459 VDD VSS PCHG WREN SEL459 BL459 BL_459 DW459 DW_459 DR459 DR_459 dido
X460 VDD VSS PCHG WREN SEL460 BL460 BL_460 DW460 DW_460 DR460 DR_460 dido
X461 VDD VSS PCHG WREN SEL461 BL461 BL_461 DW461 DW_461 DR461 DR_461 dido
X462 VDD VSS PCHG WREN SEL462 BL462 BL_462 DW462 DW_462 DR462 DR_462 dido
X463 VDD VSS PCHG WREN SEL463 BL463 BL_463 DW463 DW_463 DR463 DR_463 dido
X464 VDD VSS PCHG WREN SEL464 BL464 BL_464 DW464 DW_464 DR464 DR_464 dido
X465 VDD VSS PCHG WREN SEL465 BL465 BL_465 DW465 DW_465 DR465 DR_465 dido
X466 VDD VSS PCHG WREN SEL466 BL466 BL_466 DW466 DW_466 DR466 DR_466 dido
X467 VDD VSS PCHG WREN SEL467 BL467 BL_467 DW467 DW_467 DR467 DR_467 dido
X468 VDD VSS PCHG WREN SEL468 BL468 BL_468 DW468 DW_468 DR468 DR_468 dido
X469 VDD VSS PCHG WREN SEL469 BL469 BL_469 DW469 DW_469 DR469 DR_469 dido
X470 VDD VSS PCHG WREN SEL470 BL470 BL_470 DW470 DW_470 DR470 DR_470 dido
X471 VDD VSS PCHG WREN SEL471 BL471 BL_471 DW471 DW_471 DR471 DR_471 dido
X472 VDD VSS PCHG WREN SEL472 BL472 BL_472 DW472 DW_472 DR472 DR_472 dido
X473 VDD VSS PCHG WREN SEL473 BL473 BL_473 DW473 DW_473 DR473 DR_473 dido
X474 VDD VSS PCHG WREN SEL474 BL474 BL_474 DW474 DW_474 DR474 DR_474 dido
X475 VDD VSS PCHG WREN SEL475 BL475 BL_475 DW475 DW_475 DR475 DR_475 dido
X476 VDD VSS PCHG WREN SEL476 BL476 BL_476 DW476 DW_476 DR476 DR_476 dido
X477 VDD VSS PCHG WREN SEL477 BL477 BL_477 DW477 DW_477 DR477 DR_477 dido
X478 VDD VSS PCHG WREN SEL478 BL478 BL_478 DW478 DW_478 DR478 DR_478 dido
X479 VDD VSS PCHG WREN SEL479 BL479 BL_479 DW479 DW_479 DR479 DR_479 dido
X480 VDD VSS PCHG WREN SEL480 BL480 BL_480 DW480 DW_480 DR480 DR_480 dido
X481 VDD VSS PCHG WREN SEL481 BL481 BL_481 DW481 DW_481 DR481 DR_481 dido
X482 VDD VSS PCHG WREN SEL482 BL482 BL_482 DW482 DW_482 DR482 DR_482 dido
X483 VDD VSS PCHG WREN SEL483 BL483 BL_483 DW483 DW_483 DR483 DR_483 dido
X484 VDD VSS PCHG WREN SEL484 BL484 BL_484 DW484 DW_484 DR484 DR_484 dido
X485 VDD VSS PCHG WREN SEL485 BL485 BL_485 DW485 DW_485 DR485 DR_485 dido
X486 VDD VSS PCHG WREN SEL486 BL486 BL_486 DW486 DW_486 DR486 DR_486 dido
X487 VDD VSS PCHG WREN SEL487 BL487 BL_487 DW487 DW_487 DR487 DR_487 dido
X488 VDD VSS PCHG WREN SEL488 BL488 BL_488 DW488 DW_488 DR488 DR_488 dido
X489 VDD VSS PCHG WREN SEL489 BL489 BL_489 DW489 DW_489 DR489 DR_489 dido
X490 VDD VSS PCHG WREN SEL490 BL490 BL_490 DW490 DW_490 DR490 DR_490 dido
X491 VDD VSS PCHG WREN SEL491 BL491 BL_491 DW491 DW_491 DR491 DR_491 dido
X492 VDD VSS PCHG WREN SEL492 BL492 BL_492 DW492 DW_492 DR492 DR_492 dido
X493 VDD VSS PCHG WREN SEL493 BL493 BL_493 DW493 DW_493 DR493 DR_493 dido
X494 VDD VSS PCHG WREN SEL494 BL494 BL_494 DW494 DW_494 DR494 DR_494 dido
X495 VDD VSS PCHG WREN SEL495 BL495 BL_495 DW495 DW_495 DR495 DR_495 dido
X496 VDD VSS PCHG WREN SEL496 BL496 BL_496 DW496 DW_496 DR496 DR_496 dido
X497 VDD VSS PCHG WREN SEL497 BL497 BL_497 DW497 DW_497 DR497 DR_497 dido
X498 VDD VSS PCHG WREN SEL498 BL498 BL_498 DW498 DW_498 DR498 DR_498 dido
X499 VDD VSS PCHG WREN SEL499 BL499 BL_499 DW499 DW_499 DR499 DR_499 dido
X500 VDD VSS PCHG WREN SEL500 BL500 BL_500 DW500 DW_500 DR500 DR_500 dido
X501 VDD VSS PCHG WREN SEL501 BL501 BL_501 DW501 DW_501 DR501 DR_501 dido
X502 VDD VSS PCHG WREN SEL502 BL502 BL_502 DW502 DW_502 DR502 DR_502 dido
X503 VDD VSS PCHG WREN SEL503 BL503 BL_503 DW503 DW_503 DR503 DR_503 dido
X504 VDD VSS PCHG WREN SEL504 BL504 BL_504 DW504 DW_504 DR504 DR_504 dido
X505 VDD VSS PCHG WREN SEL505 BL505 BL_505 DW505 DW_505 DR505 DR_505 dido
X506 VDD VSS PCHG WREN SEL506 BL506 BL_506 DW506 DW_506 DR506 DR_506 dido
X507 VDD VSS PCHG WREN SEL507 BL507 BL_507 DW507 DW_507 DR507 DR_507 dido
X508 VDD VSS PCHG WREN SEL508 BL508 BL_508 DW508 DW_508 DR508 DR_508 dido
X509 VDD VSS PCHG WREN SEL509 BL509 BL_509 DW509 DW_509 DR509 DR_509 dido
X510 VDD VSS PCHG WREN SEL510 BL510 BL_510 DW510 DW_510 DR510 DR_510 dido
X511 VDD VSS PCHG WREN SEL511 BL511 BL_511 DW511 DW_511 DR511 DR_511 dido
.ends dido_arr_512

.subckt write_driver VDD VSS WREN Din DW DW_
X0 en_ WREN VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 en_ WREN VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X4 d_ Din VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X5 d_ Din VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X6 net1 Din VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X7 DW_ en_ net1 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X8 DW_ WREN net2 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
X9 net2 Din VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
X10 net3 d_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X11 DW en_ net3 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X12 DW WREN net4 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
X13 net4 d_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
.ends write_driver

.subckt del10 VDD VSS A B
X0 VDD VSS A net1 notdel
X1 VDD VSS net1 net2 notdel
X2 VDD VSS net2 net3 notdel
X3 VDD VSS net3 net4 notdel
X4 VDD VSS net4 net5 notdel
X5 VDD VSS net5 net6 notdel
X6 VDD VSS net6 net7 notdel
X7 VDD VSS net7 net8 notdel
X8 VDD VSS net8 net9 notdel
X9 VDD VSS net9 net10 notdel
X10 VDD VSS net10 net11 notdel
X11 VDD VSS A net11 net12 nand2
X12 VDD VSS net12 B not
.ends del10

.subckt ctrl VDD VSS clk cs write DBL DBL_ WREN PCHG WLEN SAEN
X0 clk_ clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 clk_ clk VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X2 WLENP clk_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 WLENP clk_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X4 VDD VSS write WREN_ not
X8 PCHG clk_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X9 PCHG clk_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
X10 DBL_ PCHG VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X11 DBL PCHG DBL_ VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X12 DBL PCHG VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X13 VDD VSS cs WLENP WLENPP nand2
X21 WLEN WLENPP VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X22 WLEN WLENPP VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
X15 VDD VSS DBL_ RBL not
X16 VDD VSS WLEN RBL SAEN_ nand2
X17 SAEN SAEN_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X18 SAEN SAEN_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
X19 WREN WREN_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X20 WREN WREN_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
.ends ctrl

.subckt input_reg8 VDD VSS clk D0 D1 D2 D3 D4 D5 D6 D7 Q0 Q1 Q2 Q3 Q4 Q5 Q6 Q7
X0 VDD VSS clk D0 Q0 in_reg
X1 VDD VSS clk D1 Q1 in_reg
X2 VDD VSS clk D2 Q2 in_reg
X3 VDD VSS clk D3 Q3 in_reg
X4 VDD VSS clk D4 Q4 in_reg
X5 VDD VSS clk D5 Q5 in_reg
X6 VDD VSS clk D6 Q6 in_reg
X7 VDD VSS clk D7 Q7 in_reg
.ends input_reg8

.subckt datain_reg128 VDD VSS clk WREN din0 din1 din2 din3 din4 din5 din6 din7 din8 din9 din10 din11 din12 din13 din14 din15 din16 din17 din18 din19 din20 din21 din22 din23 din24 din25 din26 din27 din28 din29 din30 din31 din32 din33 din34 din35 din36 din37 din38 din39 din40 din41 din42 din43 din44 din45 din46 din47 din48 din49 din50 din51 din52 din53 din54 din55 din56 din57 din58 din59 din60 din61 din62 din63 din64 din65 din66 din67 din68 din69 din70 din71 din72 din73 din74 din75 din76 din77 din78 din79 din80 din81 din82 din83 din84 din85 din86 din87 din88 din89 din90 din91 din92 din93 din94 din95 din96 din97 din98 din99 din100 din101 din102 din103 din104 din105 din106 din107 din108 din109 din110 din111 din112 din113 din114 din115 din116 din117 din118 din119 din120 din121 din122 din123 din124 din125 din126 din127 DW0 DW_0 DW1 DW_1 DW2 DW_2 DW3 DW_3 DW4 DW_4 DW5 DW_5 DW6 DW_6 DW7 DW_7 DW8 DW_8 DW9 DW_9 DW10 DW_10 DW11 DW_11 DW12 DW_12 DW13 DW_13 DW14 DW_14 DW15 DW_15 DW16 DW_16 DW17 DW_17 DW18 DW_18 DW19 DW_19 DW20 DW_20 DW21 DW_21 DW22 DW_22 DW23 DW_23 DW24 DW_24 DW25 DW_25 DW26 DW_26 DW27 DW_27 DW28 DW_28 DW29 DW_29 DW30 DW_30 DW31 DW_31 DW32 DW_32 DW33 DW_33 DW34 DW_34 DW35 DW_35 DW36 DW_36 DW37 DW_37 DW38 DW_38 DW39 DW_39 DW40 DW_40 DW41 DW_41 DW42 DW_42 DW43 DW_43 DW44 DW_44 DW45 DW_45 DW46 DW_46 DW47 DW_47 DW48 DW_48 DW49 DW_49 DW50 DW_50 DW51 DW_51 DW52 DW_52 DW53 DW_53 DW54 DW_54 DW55 DW_55 DW56 DW_56 DW57 DW_57 DW58 DW_58 DW59 DW_59 DW60 DW_60 DW61 DW_61 DW62 DW_62 DW63 DW_63 DW64 DW_64 DW65 DW_65 DW66 DW_66 DW67 DW_67 DW68 DW_68 DW69 DW_69 DW70 DW_70 DW71 DW_71 DW72 DW_72 DW73 DW_73 DW74 DW_74 DW75 DW_75 DW76 DW_76 DW77 DW_77 DW78 DW_78 DW79 DW_79 DW80 DW_80 DW81 DW_81 DW82 DW_82 DW83 DW_83 DW84 DW_84 DW85 DW_85 DW86 DW_86 DW87 DW_87 DW88 DW_88 DW89 DW_89 DW90 DW_90 DW91 DW_91 DW92 DW_92 DW93 DW_93 DW94 DW_94 DW95 DW_95 DW96 DW_96 DW97 DW_97 DW98 DW_98 DW99 DW_99 DW100 DW_100 DW101 DW_101 DW102 DW_102 DW103 DW_103 DW104 DW_104 DW105 DW_105 DW106 DW_106 DW107 DW_107 DW108 DW_108 DW109 DW_109 DW110 DW_110 DW111 DW_111 DW112 DW_112 DW113 DW_113 DW114 DW_114 DW115 DW_115 DW116 DW_116 DW117 DW_117 DW118 DW_118 DW119 DW_119 DW120 DW_120 DW121 DW_121 DW122 DW_122 DW123 DW_123 DW124 DW_124 DW125 DW_125 DW126 DW_126 DW127 DW_127
X0 VDD VSS clk din0 din_r0 in_reg
X1 VDD VSS clk din1 din_r1 in_reg
X2 VDD VSS clk din2 din_r2 in_reg
X3 VDD VSS clk din3 din_r3 in_reg
X4 VDD VSS clk din4 din_r4 in_reg
X5 VDD VSS clk din5 din_r5 in_reg
X6 VDD VSS clk din6 din_r6 in_reg
X7 VDD VSS clk din7 din_r7 in_reg
X8 VDD VSS clk din8 din_r8 in_reg
X9 VDD VSS clk din9 din_r9 in_reg
X10 VDD VSS clk din10 din_r10 in_reg
X11 VDD VSS clk din11 din_r11 in_reg
X12 VDD VSS clk din12 din_r12 in_reg
X13 VDD VSS clk din13 din_r13 in_reg
X14 VDD VSS clk din14 din_r14 in_reg
X15 VDD VSS clk din15 din_r15 in_reg
X16 VDD VSS clk din16 din_r16 in_reg
X17 VDD VSS clk din17 din_r17 in_reg
X18 VDD VSS clk din18 din_r18 in_reg
X19 VDD VSS clk din19 din_r19 in_reg
X20 VDD VSS clk din20 din_r20 in_reg
X21 VDD VSS clk din21 din_r21 in_reg
X22 VDD VSS clk din22 din_r22 in_reg
X23 VDD VSS clk din23 din_r23 in_reg
X24 VDD VSS clk din24 din_r24 in_reg
X25 VDD VSS clk din25 din_r25 in_reg
X26 VDD VSS clk din26 din_r26 in_reg
X27 VDD VSS clk din27 din_r27 in_reg
X28 VDD VSS clk din28 din_r28 in_reg
X29 VDD VSS clk din29 din_r29 in_reg
X30 VDD VSS clk din30 din_r30 in_reg
X31 VDD VSS clk din31 din_r31 in_reg
X32 VDD VSS clk din32 din_r32 in_reg
X33 VDD VSS clk din33 din_r33 in_reg
X34 VDD VSS clk din34 din_r34 in_reg
X35 VDD VSS clk din35 din_r35 in_reg
X36 VDD VSS clk din36 din_r36 in_reg
X37 VDD VSS clk din37 din_r37 in_reg
X38 VDD VSS clk din38 din_r38 in_reg
X39 VDD VSS clk din39 din_r39 in_reg
X40 VDD VSS clk din40 din_r40 in_reg
X41 VDD VSS clk din41 din_r41 in_reg
X42 VDD VSS clk din42 din_r42 in_reg
X43 VDD VSS clk din43 din_r43 in_reg
X44 VDD VSS clk din44 din_r44 in_reg
X45 VDD VSS clk din45 din_r45 in_reg
X46 VDD VSS clk din46 din_r46 in_reg
X47 VDD VSS clk din47 din_r47 in_reg
X48 VDD VSS clk din48 din_r48 in_reg
X49 VDD VSS clk din49 din_r49 in_reg
X50 VDD VSS clk din50 din_r50 in_reg
X51 VDD VSS clk din51 din_r51 in_reg
X52 VDD VSS clk din52 din_r52 in_reg
X53 VDD VSS clk din53 din_r53 in_reg
X54 VDD VSS clk din54 din_r54 in_reg
X55 VDD VSS clk din55 din_r55 in_reg
X56 VDD VSS clk din56 din_r56 in_reg
X57 VDD VSS clk din57 din_r57 in_reg
X58 VDD VSS clk din58 din_r58 in_reg
X59 VDD VSS clk din59 din_r59 in_reg
X60 VDD VSS clk din60 din_r60 in_reg
X61 VDD VSS clk din61 din_r61 in_reg
X62 VDD VSS clk din62 din_r62 in_reg
X63 VDD VSS clk din63 din_r63 in_reg
X64 VDD VSS clk din64 din_r64 in_reg
X65 VDD VSS clk din65 din_r65 in_reg
X66 VDD VSS clk din66 din_r66 in_reg
X67 VDD VSS clk din67 din_r67 in_reg
X68 VDD VSS clk din68 din_r68 in_reg
X69 VDD VSS clk din69 din_r69 in_reg
X70 VDD VSS clk din70 din_r70 in_reg
X71 VDD VSS clk din71 din_r71 in_reg
X72 VDD VSS clk din72 din_r72 in_reg
X73 VDD VSS clk din73 din_r73 in_reg
X74 VDD VSS clk din74 din_r74 in_reg
X75 VDD VSS clk din75 din_r75 in_reg
X76 VDD VSS clk din76 din_r76 in_reg
X77 VDD VSS clk din77 din_r77 in_reg
X78 VDD VSS clk din78 din_r78 in_reg
X79 VDD VSS clk din79 din_r79 in_reg
X80 VDD VSS clk din80 din_r80 in_reg
X81 VDD VSS clk din81 din_r81 in_reg
X82 VDD VSS clk din82 din_r82 in_reg
X83 VDD VSS clk din83 din_r83 in_reg
X84 VDD VSS clk din84 din_r84 in_reg
X85 VDD VSS clk din85 din_r85 in_reg
X86 VDD VSS clk din86 din_r86 in_reg
X87 VDD VSS clk din87 din_r87 in_reg
X88 VDD VSS clk din88 din_r88 in_reg
X89 VDD VSS clk din89 din_r89 in_reg
X90 VDD VSS clk din90 din_r90 in_reg
X91 VDD VSS clk din91 din_r91 in_reg
X92 VDD VSS clk din92 din_r92 in_reg
X93 VDD VSS clk din93 din_r93 in_reg
X94 VDD VSS clk din94 din_r94 in_reg
X95 VDD VSS clk din95 din_r95 in_reg
X96 VDD VSS clk din96 din_r96 in_reg
X97 VDD VSS clk din97 din_r97 in_reg
X98 VDD VSS clk din98 din_r98 in_reg
X99 VDD VSS clk din99 din_r99 in_reg
X100 VDD VSS clk din100 din_r100 in_reg
X101 VDD VSS clk din101 din_r101 in_reg
X102 VDD VSS clk din102 din_r102 in_reg
X103 VDD VSS clk din103 din_r103 in_reg
X104 VDD VSS clk din104 din_r104 in_reg
X105 VDD VSS clk din105 din_r105 in_reg
X106 VDD VSS clk din106 din_r106 in_reg
X107 VDD VSS clk din107 din_r107 in_reg
X108 VDD VSS clk din108 din_r108 in_reg
X109 VDD VSS clk din109 din_r109 in_reg
X110 VDD VSS clk din110 din_r110 in_reg
X111 VDD VSS clk din111 din_r111 in_reg
X112 VDD VSS clk din112 din_r112 in_reg
X113 VDD VSS clk din113 din_r113 in_reg
X114 VDD VSS clk din114 din_r114 in_reg
X115 VDD VSS clk din115 din_r115 in_reg
X116 VDD VSS clk din116 din_r116 in_reg
X117 VDD VSS clk din117 din_r117 in_reg
X118 VDD VSS clk din118 din_r118 in_reg
X119 VDD VSS clk din119 din_r119 in_reg
X120 VDD VSS clk din120 din_r120 in_reg
X121 VDD VSS clk din121 din_r121 in_reg
X122 VDD VSS clk din122 din_r122 in_reg
X123 VDD VSS clk din123 din_r123 in_reg
X124 VDD VSS clk din124 din_r124 in_reg
X125 VDD VSS clk din125 din_r125 in_reg
X126 VDD VSS clk din126 din_r126 in_reg
X127 VDD VSS clk din127 din_r127 in_reg
X128 VDD VSS WREN din_r0 DW0 DW_0 write_driver
X132 VDD VSS WREN din_r1 DW1 DW_1 write_driver
X136 VDD VSS WREN din_r2 DW2 DW_2 write_driver
X140 VDD VSS WREN din_r3 DW3 DW_3 write_driver
X144 VDD VSS WREN din_r4 DW4 DW_4 write_driver
X148 VDD VSS WREN din_r5 DW5 DW_5 write_driver
X152 VDD VSS WREN din_r6 DW6 DW_6 write_driver
X156 VDD VSS WREN din_r7 DW7 DW_7 write_driver
X160 VDD VSS WREN din_r8 DW8 DW_8 write_driver
X164 VDD VSS WREN din_r9 DW9 DW_9 write_driver
X168 VDD VSS WREN din_r10 DW10 DW_10 write_driver
X172 VDD VSS WREN din_r11 DW11 DW_11 write_driver
X176 VDD VSS WREN din_r12 DW12 DW_12 write_driver
X180 VDD VSS WREN din_r13 DW13 DW_13 write_driver
X184 VDD VSS WREN din_r14 DW14 DW_14 write_driver
X188 VDD VSS WREN din_r15 DW15 DW_15 write_driver
X192 VDD VSS WREN din_r16 DW16 DW_16 write_driver
X196 VDD VSS WREN din_r17 DW17 DW_17 write_driver
X200 VDD VSS WREN din_r18 DW18 DW_18 write_driver
X204 VDD VSS WREN din_r19 DW19 DW_19 write_driver
X208 VDD VSS WREN din_r20 DW20 DW_20 write_driver
X212 VDD VSS WREN din_r21 DW21 DW_21 write_driver
X216 VDD VSS WREN din_r22 DW22 DW_22 write_driver
X220 VDD VSS WREN din_r23 DW23 DW_23 write_driver
X224 VDD VSS WREN din_r24 DW24 DW_24 write_driver
X228 VDD VSS WREN din_r25 DW25 DW_25 write_driver
X232 VDD VSS WREN din_r26 DW26 DW_26 write_driver
X236 VDD VSS WREN din_r27 DW27 DW_27 write_driver
X240 VDD VSS WREN din_r28 DW28 DW_28 write_driver
X244 VDD VSS WREN din_r29 DW29 DW_29 write_driver
X248 VDD VSS WREN din_r30 DW30 DW_30 write_driver
X252 VDD VSS WREN din_r31 DW31 DW_31 write_driver
X256 VDD VSS WREN din_r32 DW32 DW_32 write_driver
X260 VDD VSS WREN din_r33 DW33 DW_33 write_driver
X264 VDD VSS WREN din_r34 DW34 DW_34 write_driver
X268 VDD VSS WREN din_r35 DW35 DW_35 write_driver
X272 VDD VSS WREN din_r36 DW36 DW_36 write_driver
X276 VDD VSS WREN din_r37 DW37 DW_37 write_driver
X280 VDD VSS WREN din_r38 DW38 DW_38 write_driver
X284 VDD VSS WREN din_r39 DW39 DW_39 write_driver
X288 VDD VSS WREN din_r40 DW40 DW_40 write_driver
X292 VDD VSS WREN din_r41 DW41 DW_41 write_driver
X296 VDD VSS WREN din_r42 DW42 DW_42 write_driver
X300 VDD VSS WREN din_r43 DW43 DW_43 write_driver
X304 VDD VSS WREN din_r44 DW44 DW_44 write_driver
X308 VDD VSS WREN din_r45 DW45 DW_45 write_driver
X312 VDD VSS WREN din_r46 DW46 DW_46 write_driver
X316 VDD VSS WREN din_r47 DW47 DW_47 write_driver
X320 VDD VSS WREN din_r48 DW48 DW_48 write_driver
X324 VDD VSS WREN din_r49 DW49 DW_49 write_driver
X328 VDD VSS WREN din_r50 DW50 DW_50 write_driver
X332 VDD VSS WREN din_r51 DW51 DW_51 write_driver
X336 VDD VSS WREN din_r52 DW52 DW_52 write_driver
X340 VDD VSS WREN din_r53 DW53 DW_53 write_driver
X344 VDD VSS WREN din_r54 DW54 DW_54 write_driver
X348 VDD VSS WREN din_r55 DW55 DW_55 write_driver
X352 VDD VSS WREN din_r56 DW56 DW_56 write_driver
X356 VDD VSS WREN din_r57 DW57 DW_57 write_driver
X360 VDD VSS WREN din_r58 DW58 DW_58 write_driver
X364 VDD VSS WREN din_r59 DW59 DW_59 write_driver
X368 VDD VSS WREN din_r60 DW60 DW_60 write_driver
X372 VDD VSS WREN din_r61 DW61 DW_61 write_driver
X376 VDD VSS WREN din_r62 DW62 DW_62 write_driver
X380 VDD VSS WREN din_r63 DW63 DW_63 write_driver
X384 VDD VSS WREN din_r64 DW64 DW_64 write_driver
X388 VDD VSS WREN din_r65 DW65 DW_65 write_driver
X392 VDD VSS WREN din_r66 DW66 DW_66 write_driver
X396 VDD VSS WREN din_r67 DW67 DW_67 write_driver
X400 VDD VSS WREN din_r68 DW68 DW_68 write_driver
X404 VDD VSS WREN din_r69 DW69 DW_69 write_driver
X408 VDD VSS WREN din_r70 DW70 DW_70 write_driver
X412 VDD VSS WREN din_r71 DW71 DW_71 write_driver
X416 VDD VSS WREN din_r72 DW72 DW_72 write_driver
X420 VDD VSS WREN din_r73 DW73 DW_73 write_driver
X424 VDD VSS WREN din_r74 DW74 DW_74 write_driver
X428 VDD VSS WREN din_r75 DW75 DW_75 write_driver
X432 VDD VSS WREN din_r76 DW76 DW_76 write_driver
X436 VDD VSS WREN din_r77 DW77 DW_77 write_driver
X440 VDD VSS WREN din_r78 DW78 DW_78 write_driver
X444 VDD VSS WREN din_r79 DW79 DW_79 write_driver
X448 VDD VSS WREN din_r80 DW80 DW_80 write_driver
X452 VDD VSS WREN din_r81 DW81 DW_81 write_driver
X456 VDD VSS WREN din_r82 DW82 DW_82 write_driver
X460 VDD VSS WREN din_r83 DW83 DW_83 write_driver
X464 VDD VSS WREN din_r84 DW84 DW_84 write_driver
X468 VDD VSS WREN din_r85 DW85 DW_85 write_driver
X472 VDD VSS WREN din_r86 DW86 DW_86 write_driver
X476 VDD VSS WREN din_r87 DW87 DW_87 write_driver
X480 VDD VSS WREN din_r88 DW88 DW_88 write_driver
X484 VDD VSS WREN din_r89 DW89 DW_89 write_driver
X488 VDD VSS WREN din_r90 DW90 DW_90 write_driver
X492 VDD VSS WREN din_r91 DW91 DW_91 write_driver
X496 VDD VSS WREN din_r92 DW92 DW_92 write_driver
X500 VDD VSS WREN din_r93 DW93 DW_93 write_driver
X504 VDD VSS WREN din_r94 DW94 DW_94 write_driver
X508 VDD VSS WREN din_r95 DW95 DW_95 write_driver
X512 VDD VSS WREN din_r96 DW96 DW_96 write_driver
X516 VDD VSS WREN din_r97 DW97 DW_97 write_driver
X520 VDD VSS WREN din_r98 DW98 DW_98 write_driver
X524 VDD VSS WREN din_r99 DW99 DW_99 write_driver
X528 VDD VSS WREN din_r100 DW100 DW_100 write_driver
X532 VDD VSS WREN din_r101 DW101 DW_101 write_driver
X536 VDD VSS WREN din_r102 DW102 DW_102 write_driver
X540 VDD VSS WREN din_r103 DW103 DW_103 write_driver
X544 VDD VSS WREN din_r104 DW104 DW_104 write_driver
X548 VDD VSS WREN din_r105 DW105 DW_105 write_driver
X552 VDD VSS WREN din_r106 DW106 DW_106 write_driver
X556 VDD VSS WREN din_r107 DW107 DW_107 write_driver
X560 VDD VSS WREN din_r108 DW108 DW_108 write_driver
X564 VDD VSS WREN din_r109 DW109 DW_109 write_driver
X568 VDD VSS WREN din_r110 DW110 DW_110 write_driver
X572 VDD VSS WREN din_r111 DW111 DW_111 write_driver
X576 VDD VSS WREN din_r112 DW112 DW_112 write_driver
X580 VDD VSS WREN din_r113 DW113 DW_113 write_driver
X584 VDD VSS WREN din_r114 DW114 DW_114 write_driver
X588 VDD VSS WREN din_r115 DW115 DW_115 write_driver
X592 VDD VSS WREN din_r116 DW116 DW_116 write_driver
X596 VDD VSS WREN din_r117 DW117 DW_117 write_driver
X600 VDD VSS WREN din_r118 DW118 DW_118 write_driver
X604 VDD VSS WREN din_r119 DW119 DW_119 write_driver
X608 VDD VSS WREN din_r120 DW120 DW_120 write_driver
X612 VDD VSS WREN din_r121 DW121 DW_121 write_driver
X616 VDD VSS WREN din_r122 DW122 DW_122 write_driver
X620 VDD VSS WREN din_r123 DW123 DW_123 write_driver
X624 VDD VSS WREN din_r124 DW124 DW_124 write_driver
X628 VDD VSS WREN din_r125 DW125 DW_125 write_driver
X632 VDD VSS WREN din_r126 DW126 DW_126 write_driver
X636 VDD VSS WREN din_r127 DW127 DW_127 write_driver
.ends datain_reg128

.subckt bit_arr_512 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL
X0 VDD VSS WL BL0 BL_0 bit_cell
X1 VDD VSS WL BL1 BL_1 bit_cell
X2 VDD VSS WL BL2 BL_2 bit_cell
X3 VDD VSS WL BL3 BL_3 bit_cell
X4 VDD VSS WL BL4 BL_4 bit_cell
X5 VDD VSS WL BL5 BL_5 bit_cell
X6 VDD VSS WL BL6 BL_6 bit_cell
X7 VDD VSS WL BL7 BL_7 bit_cell
X8 VDD VSS WL BL8 BL_8 bit_cell
X9 VDD VSS WL BL9 BL_9 bit_cell
X10 VDD VSS WL BL10 BL_10 bit_cell
X11 VDD VSS WL BL11 BL_11 bit_cell
X12 VDD VSS WL BL12 BL_12 bit_cell
X13 VDD VSS WL BL13 BL_13 bit_cell
X14 VDD VSS WL BL14 BL_14 bit_cell
X15 VDD VSS WL BL15 BL_15 bit_cell
X16 VDD VSS WL BL16 BL_16 bit_cell
X17 VDD VSS WL BL17 BL_17 bit_cell
X18 VDD VSS WL BL18 BL_18 bit_cell
X19 VDD VSS WL BL19 BL_19 bit_cell
X20 VDD VSS WL BL20 BL_20 bit_cell
X21 VDD VSS WL BL21 BL_21 bit_cell
X22 VDD VSS WL BL22 BL_22 bit_cell
X23 VDD VSS WL BL23 BL_23 bit_cell
X24 VDD VSS WL BL24 BL_24 bit_cell
X25 VDD VSS WL BL25 BL_25 bit_cell
X26 VDD VSS WL BL26 BL_26 bit_cell
X27 VDD VSS WL BL27 BL_27 bit_cell
X28 VDD VSS WL BL28 BL_28 bit_cell
X29 VDD VSS WL BL29 BL_29 bit_cell
X30 VDD VSS WL BL30 BL_30 bit_cell
X31 VDD VSS WL BL31 BL_31 bit_cell
X32 VDD VSS WL BL32 BL_32 bit_cell
X33 VDD VSS WL BL33 BL_33 bit_cell
X34 VDD VSS WL BL34 BL_34 bit_cell
X35 VDD VSS WL BL35 BL_35 bit_cell
X36 VDD VSS WL BL36 BL_36 bit_cell
X37 VDD VSS WL BL37 BL_37 bit_cell
X38 VDD VSS WL BL38 BL_38 bit_cell
X39 VDD VSS WL BL39 BL_39 bit_cell
X40 VDD VSS WL BL40 BL_40 bit_cell
X41 VDD VSS WL BL41 BL_41 bit_cell
X42 VDD VSS WL BL42 BL_42 bit_cell
X43 VDD VSS WL BL43 BL_43 bit_cell
X44 VDD VSS WL BL44 BL_44 bit_cell
X45 VDD VSS WL BL45 BL_45 bit_cell
X46 VDD VSS WL BL46 BL_46 bit_cell
X47 VDD VSS WL BL47 BL_47 bit_cell
X48 VDD VSS WL BL48 BL_48 bit_cell
X49 VDD VSS WL BL49 BL_49 bit_cell
X50 VDD VSS WL BL50 BL_50 bit_cell
X51 VDD VSS WL BL51 BL_51 bit_cell
X52 VDD VSS WL BL52 BL_52 bit_cell
X53 VDD VSS WL BL53 BL_53 bit_cell
X54 VDD VSS WL BL54 BL_54 bit_cell
X55 VDD VSS WL BL55 BL_55 bit_cell
X56 VDD VSS WL BL56 BL_56 bit_cell
X57 VDD VSS WL BL57 BL_57 bit_cell
X58 VDD VSS WL BL58 BL_58 bit_cell
X59 VDD VSS WL BL59 BL_59 bit_cell
X60 VDD VSS WL BL60 BL_60 bit_cell
X61 VDD VSS WL BL61 BL_61 bit_cell
X62 VDD VSS WL BL62 BL_62 bit_cell
X63 VDD VSS WL BL63 BL_63 bit_cell
X64 VDD VSS WL BL64 BL_64 bit_cell
X65 VDD VSS WL BL65 BL_65 bit_cell
X66 VDD VSS WL BL66 BL_66 bit_cell
X67 VDD VSS WL BL67 BL_67 bit_cell
X68 VDD VSS WL BL68 BL_68 bit_cell
X69 VDD VSS WL BL69 BL_69 bit_cell
X70 VDD VSS WL BL70 BL_70 bit_cell
X71 VDD VSS WL BL71 BL_71 bit_cell
X72 VDD VSS WL BL72 BL_72 bit_cell
X73 VDD VSS WL BL73 BL_73 bit_cell
X74 VDD VSS WL BL74 BL_74 bit_cell
X75 VDD VSS WL BL75 BL_75 bit_cell
X76 VDD VSS WL BL76 BL_76 bit_cell
X77 VDD VSS WL BL77 BL_77 bit_cell
X78 VDD VSS WL BL78 BL_78 bit_cell
X79 VDD VSS WL BL79 BL_79 bit_cell
X80 VDD VSS WL BL80 BL_80 bit_cell
X81 VDD VSS WL BL81 BL_81 bit_cell
X82 VDD VSS WL BL82 BL_82 bit_cell
X83 VDD VSS WL BL83 BL_83 bit_cell
X84 VDD VSS WL BL84 BL_84 bit_cell
X85 VDD VSS WL BL85 BL_85 bit_cell
X86 VDD VSS WL BL86 BL_86 bit_cell
X87 VDD VSS WL BL87 BL_87 bit_cell
X88 VDD VSS WL BL88 BL_88 bit_cell
X89 VDD VSS WL BL89 BL_89 bit_cell
X90 VDD VSS WL BL90 BL_90 bit_cell
X91 VDD VSS WL BL91 BL_91 bit_cell
X92 VDD VSS WL BL92 BL_92 bit_cell
X93 VDD VSS WL BL93 BL_93 bit_cell
X94 VDD VSS WL BL94 BL_94 bit_cell
X95 VDD VSS WL BL95 BL_95 bit_cell
X96 VDD VSS WL BL96 BL_96 bit_cell
X97 VDD VSS WL BL97 BL_97 bit_cell
X98 VDD VSS WL BL98 BL_98 bit_cell
X99 VDD VSS WL BL99 BL_99 bit_cell
X100 VDD VSS WL BL100 BL_100 bit_cell
X101 VDD VSS WL BL101 BL_101 bit_cell
X102 VDD VSS WL BL102 BL_102 bit_cell
X103 VDD VSS WL BL103 BL_103 bit_cell
X104 VDD VSS WL BL104 BL_104 bit_cell
X105 VDD VSS WL BL105 BL_105 bit_cell
X106 VDD VSS WL BL106 BL_106 bit_cell
X107 VDD VSS WL BL107 BL_107 bit_cell
X108 VDD VSS WL BL108 BL_108 bit_cell
X109 VDD VSS WL BL109 BL_109 bit_cell
X110 VDD VSS WL BL110 BL_110 bit_cell
X111 VDD VSS WL BL111 BL_111 bit_cell
X112 VDD VSS WL BL112 BL_112 bit_cell
X113 VDD VSS WL BL113 BL_113 bit_cell
X114 VDD VSS WL BL114 BL_114 bit_cell
X115 VDD VSS WL BL115 BL_115 bit_cell
X116 VDD VSS WL BL116 BL_116 bit_cell
X117 VDD VSS WL BL117 BL_117 bit_cell
X118 VDD VSS WL BL118 BL_118 bit_cell
X119 VDD VSS WL BL119 BL_119 bit_cell
X120 VDD VSS WL BL120 BL_120 bit_cell
X121 VDD VSS WL BL121 BL_121 bit_cell
X122 VDD VSS WL BL122 BL_122 bit_cell
X123 VDD VSS WL BL123 BL_123 bit_cell
X124 VDD VSS WL BL124 BL_124 bit_cell
X125 VDD VSS WL BL125 BL_125 bit_cell
X126 VDD VSS WL BL126 BL_126 bit_cell
X127 VDD VSS WL BL127 BL_127 bit_cell
X128 VDD VSS WL BL128 BL_128 bit_cell
X129 VDD VSS WL BL129 BL_129 bit_cell
X130 VDD VSS WL BL130 BL_130 bit_cell
X131 VDD VSS WL BL131 BL_131 bit_cell
X132 VDD VSS WL BL132 BL_132 bit_cell
X133 VDD VSS WL BL133 BL_133 bit_cell
X134 VDD VSS WL BL134 BL_134 bit_cell
X135 VDD VSS WL BL135 BL_135 bit_cell
X136 VDD VSS WL BL136 BL_136 bit_cell
X137 VDD VSS WL BL137 BL_137 bit_cell
X138 VDD VSS WL BL138 BL_138 bit_cell
X139 VDD VSS WL BL139 BL_139 bit_cell
X140 VDD VSS WL BL140 BL_140 bit_cell
X141 VDD VSS WL BL141 BL_141 bit_cell
X142 VDD VSS WL BL142 BL_142 bit_cell
X143 VDD VSS WL BL143 BL_143 bit_cell
X144 VDD VSS WL BL144 BL_144 bit_cell
X145 VDD VSS WL BL145 BL_145 bit_cell
X146 VDD VSS WL BL146 BL_146 bit_cell
X147 VDD VSS WL BL147 BL_147 bit_cell
X148 VDD VSS WL BL148 BL_148 bit_cell
X149 VDD VSS WL BL149 BL_149 bit_cell
X150 VDD VSS WL BL150 BL_150 bit_cell
X151 VDD VSS WL BL151 BL_151 bit_cell
X152 VDD VSS WL BL152 BL_152 bit_cell
X153 VDD VSS WL BL153 BL_153 bit_cell
X154 VDD VSS WL BL154 BL_154 bit_cell
X155 VDD VSS WL BL155 BL_155 bit_cell
X156 VDD VSS WL BL156 BL_156 bit_cell
X157 VDD VSS WL BL157 BL_157 bit_cell
X158 VDD VSS WL BL158 BL_158 bit_cell
X159 VDD VSS WL BL159 BL_159 bit_cell
X160 VDD VSS WL BL160 BL_160 bit_cell
X161 VDD VSS WL BL161 BL_161 bit_cell
X162 VDD VSS WL BL162 BL_162 bit_cell
X163 VDD VSS WL BL163 BL_163 bit_cell
X164 VDD VSS WL BL164 BL_164 bit_cell
X165 VDD VSS WL BL165 BL_165 bit_cell
X166 VDD VSS WL BL166 BL_166 bit_cell
X167 VDD VSS WL BL167 BL_167 bit_cell
X168 VDD VSS WL BL168 BL_168 bit_cell
X169 VDD VSS WL BL169 BL_169 bit_cell
X170 VDD VSS WL BL170 BL_170 bit_cell
X171 VDD VSS WL BL171 BL_171 bit_cell
X172 VDD VSS WL BL172 BL_172 bit_cell
X173 VDD VSS WL BL173 BL_173 bit_cell
X174 VDD VSS WL BL174 BL_174 bit_cell
X175 VDD VSS WL BL175 BL_175 bit_cell
X176 VDD VSS WL BL176 BL_176 bit_cell
X177 VDD VSS WL BL177 BL_177 bit_cell
X178 VDD VSS WL BL178 BL_178 bit_cell
X179 VDD VSS WL BL179 BL_179 bit_cell
X180 VDD VSS WL BL180 BL_180 bit_cell
X181 VDD VSS WL BL181 BL_181 bit_cell
X182 VDD VSS WL BL182 BL_182 bit_cell
X183 VDD VSS WL BL183 BL_183 bit_cell
X184 VDD VSS WL BL184 BL_184 bit_cell
X185 VDD VSS WL BL185 BL_185 bit_cell
X186 VDD VSS WL BL186 BL_186 bit_cell
X187 VDD VSS WL BL187 BL_187 bit_cell
X188 VDD VSS WL BL188 BL_188 bit_cell
X189 VDD VSS WL BL189 BL_189 bit_cell
X190 VDD VSS WL BL190 BL_190 bit_cell
X191 VDD VSS WL BL191 BL_191 bit_cell
X192 VDD VSS WL BL192 BL_192 bit_cell
X193 VDD VSS WL BL193 BL_193 bit_cell
X194 VDD VSS WL BL194 BL_194 bit_cell
X195 VDD VSS WL BL195 BL_195 bit_cell
X196 VDD VSS WL BL196 BL_196 bit_cell
X197 VDD VSS WL BL197 BL_197 bit_cell
X198 VDD VSS WL BL198 BL_198 bit_cell
X199 VDD VSS WL BL199 BL_199 bit_cell
X200 VDD VSS WL BL200 BL_200 bit_cell
X201 VDD VSS WL BL201 BL_201 bit_cell
X202 VDD VSS WL BL202 BL_202 bit_cell
X203 VDD VSS WL BL203 BL_203 bit_cell
X204 VDD VSS WL BL204 BL_204 bit_cell
X205 VDD VSS WL BL205 BL_205 bit_cell
X206 VDD VSS WL BL206 BL_206 bit_cell
X207 VDD VSS WL BL207 BL_207 bit_cell
X208 VDD VSS WL BL208 BL_208 bit_cell
X209 VDD VSS WL BL209 BL_209 bit_cell
X210 VDD VSS WL BL210 BL_210 bit_cell
X211 VDD VSS WL BL211 BL_211 bit_cell
X212 VDD VSS WL BL212 BL_212 bit_cell
X213 VDD VSS WL BL213 BL_213 bit_cell
X214 VDD VSS WL BL214 BL_214 bit_cell
X215 VDD VSS WL BL215 BL_215 bit_cell
X216 VDD VSS WL BL216 BL_216 bit_cell
X217 VDD VSS WL BL217 BL_217 bit_cell
X218 VDD VSS WL BL218 BL_218 bit_cell
X219 VDD VSS WL BL219 BL_219 bit_cell
X220 VDD VSS WL BL220 BL_220 bit_cell
X221 VDD VSS WL BL221 BL_221 bit_cell
X222 VDD VSS WL BL222 BL_222 bit_cell
X223 VDD VSS WL BL223 BL_223 bit_cell
X224 VDD VSS WL BL224 BL_224 bit_cell
X225 VDD VSS WL BL225 BL_225 bit_cell
X226 VDD VSS WL BL226 BL_226 bit_cell
X227 VDD VSS WL BL227 BL_227 bit_cell
X228 VDD VSS WL BL228 BL_228 bit_cell
X229 VDD VSS WL BL229 BL_229 bit_cell
X230 VDD VSS WL BL230 BL_230 bit_cell
X231 VDD VSS WL BL231 BL_231 bit_cell
X232 VDD VSS WL BL232 BL_232 bit_cell
X233 VDD VSS WL BL233 BL_233 bit_cell
X234 VDD VSS WL BL234 BL_234 bit_cell
X235 VDD VSS WL BL235 BL_235 bit_cell
X236 VDD VSS WL BL236 BL_236 bit_cell
X237 VDD VSS WL BL237 BL_237 bit_cell
X238 VDD VSS WL BL238 BL_238 bit_cell
X239 VDD VSS WL BL239 BL_239 bit_cell
X240 VDD VSS WL BL240 BL_240 bit_cell
X241 VDD VSS WL BL241 BL_241 bit_cell
X242 VDD VSS WL BL242 BL_242 bit_cell
X243 VDD VSS WL BL243 BL_243 bit_cell
X244 VDD VSS WL BL244 BL_244 bit_cell
X245 VDD VSS WL BL245 BL_245 bit_cell
X246 VDD VSS WL BL246 BL_246 bit_cell
X247 VDD VSS WL BL247 BL_247 bit_cell
X248 VDD VSS WL BL248 BL_248 bit_cell
X249 VDD VSS WL BL249 BL_249 bit_cell
X250 VDD VSS WL BL250 BL_250 bit_cell
X251 VDD VSS WL BL251 BL_251 bit_cell
X252 VDD VSS WL BL252 BL_252 bit_cell
X253 VDD VSS WL BL253 BL_253 bit_cell
X254 VDD VSS WL BL254 BL_254 bit_cell
X255 VDD VSS WL BL255 BL_255 bit_cell
X256 VDD VSS WL BL256 BL_256 bit_cell
X257 VDD VSS WL BL257 BL_257 bit_cell
X258 VDD VSS WL BL258 BL_258 bit_cell
X259 VDD VSS WL BL259 BL_259 bit_cell
X260 VDD VSS WL BL260 BL_260 bit_cell
X261 VDD VSS WL BL261 BL_261 bit_cell
X262 VDD VSS WL BL262 BL_262 bit_cell
X263 VDD VSS WL BL263 BL_263 bit_cell
X264 VDD VSS WL BL264 BL_264 bit_cell
X265 VDD VSS WL BL265 BL_265 bit_cell
X266 VDD VSS WL BL266 BL_266 bit_cell
X267 VDD VSS WL BL267 BL_267 bit_cell
X268 VDD VSS WL BL268 BL_268 bit_cell
X269 VDD VSS WL BL269 BL_269 bit_cell
X270 VDD VSS WL BL270 BL_270 bit_cell
X271 VDD VSS WL BL271 BL_271 bit_cell
X272 VDD VSS WL BL272 BL_272 bit_cell
X273 VDD VSS WL BL273 BL_273 bit_cell
X274 VDD VSS WL BL274 BL_274 bit_cell
X275 VDD VSS WL BL275 BL_275 bit_cell
X276 VDD VSS WL BL276 BL_276 bit_cell
X277 VDD VSS WL BL277 BL_277 bit_cell
X278 VDD VSS WL BL278 BL_278 bit_cell
X279 VDD VSS WL BL279 BL_279 bit_cell
X280 VDD VSS WL BL280 BL_280 bit_cell
X281 VDD VSS WL BL281 BL_281 bit_cell
X282 VDD VSS WL BL282 BL_282 bit_cell
X283 VDD VSS WL BL283 BL_283 bit_cell
X284 VDD VSS WL BL284 BL_284 bit_cell
X285 VDD VSS WL BL285 BL_285 bit_cell
X286 VDD VSS WL BL286 BL_286 bit_cell
X287 VDD VSS WL BL287 BL_287 bit_cell
X288 VDD VSS WL BL288 BL_288 bit_cell
X289 VDD VSS WL BL289 BL_289 bit_cell
X290 VDD VSS WL BL290 BL_290 bit_cell
X291 VDD VSS WL BL291 BL_291 bit_cell
X292 VDD VSS WL BL292 BL_292 bit_cell
X293 VDD VSS WL BL293 BL_293 bit_cell
X294 VDD VSS WL BL294 BL_294 bit_cell
X295 VDD VSS WL BL295 BL_295 bit_cell
X296 VDD VSS WL BL296 BL_296 bit_cell
X297 VDD VSS WL BL297 BL_297 bit_cell
X298 VDD VSS WL BL298 BL_298 bit_cell
X299 VDD VSS WL BL299 BL_299 bit_cell
X300 VDD VSS WL BL300 BL_300 bit_cell
X301 VDD VSS WL BL301 BL_301 bit_cell
X302 VDD VSS WL BL302 BL_302 bit_cell
X303 VDD VSS WL BL303 BL_303 bit_cell
X304 VDD VSS WL BL304 BL_304 bit_cell
X305 VDD VSS WL BL305 BL_305 bit_cell
X306 VDD VSS WL BL306 BL_306 bit_cell
X307 VDD VSS WL BL307 BL_307 bit_cell
X308 VDD VSS WL BL308 BL_308 bit_cell
X309 VDD VSS WL BL309 BL_309 bit_cell
X310 VDD VSS WL BL310 BL_310 bit_cell
X311 VDD VSS WL BL311 BL_311 bit_cell
X312 VDD VSS WL BL312 BL_312 bit_cell
X313 VDD VSS WL BL313 BL_313 bit_cell
X314 VDD VSS WL BL314 BL_314 bit_cell
X315 VDD VSS WL BL315 BL_315 bit_cell
X316 VDD VSS WL BL316 BL_316 bit_cell
X317 VDD VSS WL BL317 BL_317 bit_cell
X318 VDD VSS WL BL318 BL_318 bit_cell
X319 VDD VSS WL BL319 BL_319 bit_cell
X320 VDD VSS WL BL320 BL_320 bit_cell
X321 VDD VSS WL BL321 BL_321 bit_cell
X322 VDD VSS WL BL322 BL_322 bit_cell
X323 VDD VSS WL BL323 BL_323 bit_cell
X324 VDD VSS WL BL324 BL_324 bit_cell
X325 VDD VSS WL BL325 BL_325 bit_cell
X326 VDD VSS WL BL326 BL_326 bit_cell
X327 VDD VSS WL BL327 BL_327 bit_cell
X328 VDD VSS WL BL328 BL_328 bit_cell
X329 VDD VSS WL BL329 BL_329 bit_cell
X330 VDD VSS WL BL330 BL_330 bit_cell
X331 VDD VSS WL BL331 BL_331 bit_cell
X332 VDD VSS WL BL332 BL_332 bit_cell
X333 VDD VSS WL BL333 BL_333 bit_cell
X334 VDD VSS WL BL334 BL_334 bit_cell
X335 VDD VSS WL BL335 BL_335 bit_cell
X336 VDD VSS WL BL336 BL_336 bit_cell
X337 VDD VSS WL BL337 BL_337 bit_cell
X338 VDD VSS WL BL338 BL_338 bit_cell
X339 VDD VSS WL BL339 BL_339 bit_cell
X340 VDD VSS WL BL340 BL_340 bit_cell
X341 VDD VSS WL BL341 BL_341 bit_cell
X342 VDD VSS WL BL342 BL_342 bit_cell
X343 VDD VSS WL BL343 BL_343 bit_cell
X344 VDD VSS WL BL344 BL_344 bit_cell
X345 VDD VSS WL BL345 BL_345 bit_cell
X346 VDD VSS WL BL346 BL_346 bit_cell
X347 VDD VSS WL BL347 BL_347 bit_cell
X348 VDD VSS WL BL348 BL_348 bit_cell
X349 VDD VSS WL BL349 BL_349 bit_cell
X350 VDD VSS WL BL350 BL_350 bit_cell
X351 VDD VSS WL BL351 BL_351 bit_cell
X352 VDD VSS WL BL352 BL_352 bit_cell
X353 VDD VSS WL BL353 BL_353 bit_cell
X354 VDD VSS WL BL354 BL_354 bit_cell
X355 VDD VSS WL BL355 BL_355 bit_cell
X356 VDD VSS WL BL356 BL_356 bit_cell
X357 VDD VSS WL BL357 BL_357 bit_cell
X358 VDD VSS WL BL358 BL_358 bit_cell
X359 VDD VSS WL BL359 BL_359 bit_cell
X360 VDD VSS WL BL360 BL_360 bit_cell
X361 VDD VSS WL BL361 BL_361 bit_cell
X362 VDD VSS WL BL362 BL_362 bit_cell
X363 VDD VSS WL BL363 BL_363 bit_cell
X364 VDD VSS WL BL364 BL_364 bit_cell
X365 VDD VSS WL BL365 BL_365 bit_cell
X366 VDD VSS WL BL366 BL_366 bit_cell
X367 VDD VSS WL BL367 BL_367 bit_cell
X368 VDD VSS WL BL368 BL_368 bit_cell
X369 VDD VSS WL BL369 BL_369 bit_cell
X370 VDD VSS WL BL370 BL_370 bit_cell
X371 VDD VSS WL BL371 BL_371 bit_cell
X372 VDD VSS WL BL372 BL_372 bit_cell
X373 VDD VSS WL BL373 BL_373 bit_cell
X374 VDD VSS WL BL374 BL_374 bit_cell
X375 VDD VSS WL BL375 BL_375 bit_cell
X376 VDD VSS WL BL376 BL_376 bit_cell
X377 VDD VSS WL BL377 BL_377 bit_cell
X378 VDD VSS WL BL378 BL_378 bit_cell
X379 VDD VSS WL BL379 BL_379 bit_cell
X380 VDD VSS WL BL380 BL_380 bit_cell
X381 VDD VSS WL BL381 BL_381 bit_cell
X382 VDD VSS WL BL382 BL_382 bit_cell
X383 VDD VSS WL BL383 BL_383 bit_cell
X384 VDD VSS WL BL384 BL_384 bit_cell
X385 VDD VSS WL BL385 BL_385 bit_cell
X386 VDD VSS WL BL386 BL_386 bit_cell
X387 VDD VSS WL BL387 BL_387 bit_cell
X388 VDD VSS WL BL388 BL_388 bit_cell
X389 VDD VSS WL BL389 BL_389 bit_cell
X390 VDD VSS WL BL390 BL_390 bit_cell
X391 VDD VSS WL BL391 BL_391 bit_cell
X392 VDD VSS WL BL392 BL_392 bit_cell
X393 VDD VSS WL BL393 BL_393 bit_cell
X394 VDD VSS WL BL394 BL_394 bit_cell
X395 VDD VSS WL BL395 BL_395 bit_cell
X396 VDD VSS WL BL396 BL_396 bit_cell
X397 VDD VSS WL BL397 BL_397 bit_cell
X398 VDD VSS WL BL398 BL_398 bit_cell
X399 VDD VSS WL BL399 BL_399 bit_cell
X400 VDD VSS WL BL400 BL_400 bit_cell
X401 VDD VSS WL BL401 BL_401 bit_cell
X402 VDD VSS WL BL402 BL_402 bit_cell
X403 VDD VSS WL BL403 BL_403 bit_cell
X404 VDD VSS WL BL404 BL_404 bit_cell
X405 VDD VSS WL BL405 BL_405 bit_cell
X406 VDD VSS WL BL406 BL_406 bit_cell
X407 VDD VSS WL BL407 BL_407 bit_cell
X408 VDD VSS WL BL408 BL_408 bit_cell
X409 VDD VSS WL BL409 BL_409 bit_cell
X410 VDD VSS WL BL410 BL_410 bit_cell
X411 VDD VSS WL BL411 BL_411 bit_cell
X412 VDD VSS WL BL412 BL_412 bit_cell
X413 VDD VSS WL BL413 BL_413 bit_cell
X414 VDD VSS WL BL414 BL_414 bit_cell
X415 VDD VSS WL BL415 BL_415 bit_cell
X416 VDD VSS WL BL416 BL_416 bit_cell
X417 VDD VSS WL BL417 BL_417 bit_cell
X418 VDD VSS WL BL418 BL_418 bit_cell
X419 VDD VSS WL BL419 BL_419 bit_cell
X420 VDD VSS WL BL420 BL_420 bit_cell
X421 VDD VSS WL BL421 BL_421 bit_cell
X422 VDD VSS WL BL422 BL_422 bit_cell
X423 VDD VSS WL BL423 BL_423 bit_cell
X424 VDD VSS WL BL424 BL_424 bit_cell
X425 VDD VSS WL BL425 BL_425 bit_cell
X426 VDD VSS WL BL426 BL_426 bit_cell
X427 VDD VSS WL BL427 BL_427 bit_cell
X428 VDD VSS WL BL428 BL_428 bit_cell
X429 VDD VSS WL BL429 BL_429 bit_cell
X430 VDD VSS WL BL430 BL_430 bit_cell
X431 VDD VSS WL BL431 BL_431 bit_cell
X432 VDD VSS WL BL432 BL_432 bit_cell
X433 VDD VSS WL BL433 BL_433 bit_cell
X434 VDD VSS WL BL434 BL_434 bit_cell
X435 VDD VSS WL BL435 BL_435 bit_cell
X436 VDD VSS WL BL436 BL_436 bit_cell
X437 VDD VSS WL BL437 BL_437 bit_cell
X438 VDD VSS WL BL438 BL_438 bit_cell
X439 VDD VSS WL BL439 BL_439 bit_cell
X440 VDD VSS WL BL440 BL_440 bit_cell
X441 VDD VSS WL BL441 BL_441 bit_cell
X442 VDD VSS WL BL442 BL_442 bit_cell
X443 VDD VSS WL BL443 BL_443 bit_cell
X444 VDD VSS WL BL444 BL_444 bit_cell
X445 VDD VSS WL BL445 BL_445 bit_cell
X446 VDD VSS WL BL446 BL_446 bit_cell
X447 VDD VSS WL BL447 BL_447 bit_cell
X448 VDD VSS WL BL448 BL_448 bit_cell
X449 VDD VSS WL BL449 BL_449 bit_cell
X450 VDD VSS WL BL450 BL_450 bit_cell
X451 VDD VSS WL BL451 BL_451 bit_cell
X452 VDD VSS WL BL452 BL_452 bit_cell
X453 VDD VSS WL BL453 BL_453 bit_cell
X454 VDD VSS WL BL454 BL_454 bit_cell
X455 VDD VSS WL BL455 BL_455 bit_cell
X456 VDD VSS WL BL456 BL_456 bit_cell
X457 VDD VSS WL BL457 BL_457 bit_cell
X458 VDD VSS WL BL458 BL_458 bit_cell
X459 VDD VSS WL BL459 BL_459 bit_cell
X460 VDD VSS WL BL460 BL_460 bit_cell
X461 VDD VSS WL BL461 BL_461 bit_cell
X462 VDD VSS WL BL462 BL_462 bit_cell
X463 VDD VSS WL BL463 BL_463 bit_cell
X464 VDD VSS WL BL464 BL_464 bit_cell
X465 VDD VSS WL BL465 BL_465 bit_cell
X466 VDD VSS WL BL466 BL_466 bit_cell
X467 VDD VSS WL BL467 BL_467 bit_cell
X468 VDD VSS WL BL468 BL_468 bit_cell
X469 VDD VSS WL BL469 BL_469 bit_cell
X470 VDD VSS WL BL470 BL_470 bit_cell
X471 VDD VSS WL BL471 BL_471 bit_cell
X472 VDD VSS WL BL472 BL_472 bit_cell
X473 VDD VSS WL BL473 BL_473 bit_cell
X474 VDD VSS WL BL474 BL_474 bit_cell
X475 VDD VSS WL BL475 BL_475 bit_cell
X476 VDD VSS WL BL476 BL_476 bit_cell
X477 VDD VSS WL BL477 BL_477 bit_cell
X478 VDD VSS WL BL478 BL_478 bit_cell
X479 VDD VSS WL BL479 BL_479 bit_cell
X480 VDD VSS WL BL480 BL_480 bit_cell
X481 VDD VSS WL BL481 BL_481 bit_cell
X482 VDD VSS WL BL482 BL_482 bit_cell
X483 VDD VSS WL BL483 BL_483 bit_cell
X484 VDD VSS WL BL484 BL_484 bit_cell
X485 VDD VSS WL BL485 BL_485 bit_cell
X486 VDD VSS WL BL486 BL_486 bit_cell
X487 VDD VSS WL BL487 BL_487 bit_cell
X488 VDD VSS WL BL488 BL_488 bit_cell
X489 VDD VSS WL BL489 BL_489 bit_cell
X490 VDD VSS WL BL490 BL_490 bit_cell
X491 VDD VSS WL BL491 BL_491 bit_cell
X492 VDD VSS WL BL492 BL_492 bit_cell
X493 VDD VSS WL BL493 BL_493 bit_cell
X494 VDD VSS WL BL494 BL_494 bit_cell
X495 VDD VSS WL BL495 BL_495 bit_cell
X496 VDD VSS WL BL496 BL_496 bit_cell
X497 VDD VSS WL BL497 BL_497 bit_cell
X498 VDD VSS WL BL498 BL_498 bit_cell
X499 VDD VSS WL BL499 BL_499 bit_cell
X500 VDD VSS WL BL500 BL_500 bit_cell
X501 VDD VSS WL BL501 BL_501 bit_cell
X502 VDD VSS WL BL502 BL_502 bit_cell
X503 VDD VSS WL BL503 BL_503 bit_cell
X504 VDD VSS WL BL504 BL_504 bit_cell
X505 VDD VSS WL BL505 BL_505 bit_cell
X506 VDD VSS WL BL506 BL_506 bit_cell
X507 VDD VSS WL BL507 BL_507 bit_cell
X508 VDD VSS WL BL508 BL_508 bit_cell
X509 VDD VSS WL BL509 BL_509 bit_cell
X510 VDD VSS WL BL510 BL_510 bit_cell
X511 VDD VSS WL BL511 BL_511 bit_cell
.ends bit_arr_512

.subckt dmy_arr_32 VDD VSS WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 DBL DBL_
X0 VDD VSS WL0 DBL DBL_ dmy_cell
X1 VDD VSS WL1 DBL DBL_ dmy_cell
X2 VDD VSS WL2 DBL DBL_ dmy_cell
X3 VDD VSS WL3 DBL DBL_ dmy_cell
X4 VDD VSS WL4 DBL DBL_ dmy_cell
X5 VDD VSS WL5 DBL DBL_ dmy_cell
X6 VDD VSS WL6 DBL DBL_ dmy_cell
X7 VDD VSS WL7 DBL DBL_ dmy_cell
X8 VDD VSS WL8 DBL DBL_ dmy_cell
X9 VDD VSS WL9 DBL DBL_ dmy_cell
X10 VDD VSS WL10 DBL DBL_ dmy_cell
X11 VDD VSS WL11 DBL DBL_ dmy_cell
X12 VDD VSS WL12 DBL DBL_ dmy_cell
X13 VDD VSS WL13 DBL DBL_ dmy_cell
X14 VDD VSS WL14 DBL DBL_ dmy_cell
X15 VDD VSS WL15 DBL DBL_ dmy_cell
X16 VDD VSS WL16 DBL DBL_ dmy_cell
X17 VDD VSS WL17 DBL DBL_ dmy_cell
X18 VDD VSS WL18 DBL DBL_ dmy_cell
X19 VDD VSS WL19 DBL DBL_ dmy_cell
X20 VDD VSS WL20 DBL DBL_ dmy_cell
X21 VDD VSS WL21 DBL DBL_ dmy_cell
X22 VDD VSS WL22 DBL DBL_ dmy_cell
X23 VDD VSS WL23 DBL DBL_ dmy_cell
X24 VDD VSS WL24 DBL DBL_ dmy_cell
X25 VDD VSS WL25 DBL DBL_ dmy_cell
X26 VDD VSS WL26 DBL DBL_ dmy_cell
X27 VDD VSS WL27 DBL DBL_ dmy_cell
X28 VDD VSS WL28 DBL DBL_ dmy_cell
X29 VDD VSS WL29 DBL DBL_ dmy_cell
X30 VDD VSS WL30 DBL DBL_ dmy_cell
X31 VDD VSS WL31 DBL DBL_ dmy_cell
.ends dmy_arr_32

.subckt se_arr_128 VDD VSS SAEN BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 SB0 SB1 SB2 SB3 SB4 SB5 SB6 SB7 SB8 SB9 SB10 SB11 SB12 SB13 SB14 SB15 SB16 SB17 SB18 SB19 SB20 SB21 SB22 SB23 SB24 SB25 SB26 SB27 SB28 SB29 SB30 SB31 SB32 SB33 SB34 SB35 SB36 SB37 SB38 SB39 SB40 SB41 SB42 SB43 SB44 SB45 SB46 SB47 SB48 SB49 SB50 SB51 SB52 SB53 SB54 SB55 SB56 SB57 SB58 SB59 SB60 SB61 SB62 SB63 SB64 SB65 SB66 SB67 SB68 SB69 SB70 SB71 SB72 SB73 SB74 SB75 SB76 SB77 SB78 SB79 SB80 SB81 SB82 SB83 SB84 SB85 SB86 SB87 SB88 SB89 SB90 SB91 SB92 SB93 SB94 SB95 SB96 SB97 SB98 SB99 SB100 SB101 SB102 SB103 SB104 SB105 SB106 SB107 SB108 SB109 SB110 SB111 SB112 SB113 SB114 SB115 SB116 SB117 SB118 SB119 SB120 SB121 SB122 SB123 SB124 SB125 SB126 SB127
X0 VDD VSS SAEN BL0 BL_0 SB0 se_cell
X1 VDD VSS SAEN BL1 BL_1 SB1 se_cell
X2 VDD VSS SAEN BL2 BL_2 SB2 se_cell
X3 VDD VSS SAEN BL3 BL_3 SB3 se_cell
X4 VDD VSS SAEN BL4 BL_4 SB4 se_cell
X5 VDD VSS SAEN BL5 BL_5 SB5 se_cell
X6 VDD VSS SAEN BL6 BL_6 SB6 se_cell
X7 VDD VSS SAEN BL7 BL_7 SB7 se_cell
X8 VDD VSS SAEN BL8 BL_8 SB8 se_cell
X9 VDD VSS SAEN BL9 BL_9 SB9 se_cell
X10 VDD VSS SAEN BL10 BL_10 SB10 se_cell
X11 VDD VSS SAEN BL11 BL_11 SB11 se_cell
X12 VDD VSS SAEN BL12 BL_12 SB12 se_cell
X13 VDD VSS SAEN BL13 BL_13 SB13 se_cell
X14 VDD VSS SAEN BL14 BL_14 SB14 se_cell
X15 VDD VSS SAEN BL15 BL_15 SB15 se_cell
X16 VDD VSS SAEN BL16 BL_16 SB16 se_cell
X17 VDD VSS SAEN BL17 BL_17 SB17 se_cell
X18 VDD VSS SAEN BL18 BL_18 SB18 se_cell
X19 VDD VSS SAEN BL19 BL_19 SB19 se_cell
X20 VDD VSS SAEN BL20 BL_20 SB20 se_cell
X21 VDD VSS SAEN BL21 BL_21 SB21 se_cell
X22 VDD VSS SAEN BL22 BL_22 SB22 se_cell
X23 VDD VSS SAEN BL23 BL_23 SB23 se_cell
X24 VDD VSS SAEN BL24 BL_24 SB24 se_cell
X25 VDD VSS SAEN BL25 BL_25 SB25 se_cell
X26 VDD VSS SAEN BL26 BL_26 SB26 se_cell
X27 VDD VSS SAEN BL27 BL_27 SB27 se_cell
X28 VDD VSS SAEN BL28 BL_28 SB28 se_cell
X29 VDD VSS SAEN BL29 BL_29 SB29 se_cell
X30 VDD VSS SAEN BL30 BL_30 SB30 se_cell
X31 VDD VSS SAEN BL31 BL_31 SB31 se_cell
X32 VDD VSS SAEN BL32 BL_32 SB32 se_cell
X33 VDD VSS SAEN BL33 BL_33 SB33 se_cell
X34 VDD VSS SAEN BL34 BL_34 SB34 se_cell
X35 VDD VSS SAEN BL35 BL_35 SB35 se_cell
X36 VDD VSS SAEN BL36 BL_36 SB36 se_cell
X37 VDD VSS SAEN BL37 BL_37 SB37 se_cell
X38 VDD VSS SAEN BL38 BL_38 SB38 se_cell
X39 VDD VSS SAEN BL39 BL_39 SB39 se_cell
X40 VDD VSS SAEN BL40 BL_40 SB40 se_cell
X41 VDD VSS SAEN BL41 BL_41 SB41 se_cell
X42 VDD VSS SAEN BL42 BL_42 SB42 se_cell
X43 VDD VSS SAEN BL43 BL_43 SB43 se_cell
X44 VDD VSS SAEN BL44 BL_44 SB44 se_cell
X45 VDD VSS SAEN BL45 BL_45 SB45 se_cell
X46 VDD VSS SAEN BL46 BL_46 SB46 se_cell
X47 VDD VSS SAEN BL47 BL_47 SB47 se_cell
X48 VDD VSS SAEN BL48 BL_48 SB48 se_cell
X49 VDD VSS SAEN BL49 BL_49 SB49 se_cell
X50 VDD VSS SAEN BL50 BL_50 SB50 se_cell
X51 VDD VSS SAEN BL51 BL_51 SB51 se_cell
X52 VDD VSS SAEN BL52 BL_52 SB52 se_cell
X53 VDD VSS SAEN BL53 BL_53 SB53 se_cell
X54 VDD VSS SAEN BL54 BL_54 SB54 se_cell
X55 VDD VSS SAEN BL55 BL_55 SB55 se_cell
X56 VDD VSS SAEN BL56 BL_56 SB56 se_cell
X57 VDD VSS SAEN BL57 BL_57 SB57 se_cell
X58 VDD VSS SAEN BL58 BL_58 SB58 se_cell
X59 VDD VSS SAEN BL59 BL_59 SB59 se_cell
X60 VDD VSS SAEN BL60 BL_60 SB60 se_cell
X61 VDD VSS SAEN BL61 BL_61 SB61 se_cell
X62 VDD VSS SAEN BL62 BL_62 SB62 se_cell
X63 VDD VSS SAEN BL63 BL_63 SB63 se_cell
X64 VDD VSS SAEN BL64 BL_64 SB64 se_cell
X65 VDD VSS SAEN BL65 BL_65 SB65 se_cell
X66 VDD VSS SAEN BL66 BL_66 SB66 se_cell
X67 VDD VSS SAEN BL67 BL_67 SB67 se_cell
X68 VDD VSS SAEN BL68 BL_68 SB68 se_cell
X69 VDD VSS SAEN BL69 BL_69 SB69 se_cell
X70 VDD VSS SAEN BL70 BL_70 SB70 se_cell
X71 VDD VSS SAEN BL71 BL_71 SB71 se_cell
X72 VDD VSS SAEN BL72 BL_72 SB72 se_cell
X73 VDD VSS SAEN BL73 BL_73 SB73 se_cell
X74 VDD VSS SAEN BL74 BL_74 SB74 se_cell
X75 VDD VSS SAEN BL75 BL_75 SB75 se_cell
X76 VDD VSS SAEN BL76 BL_76 SB76 se_cell
X77 VDD VSS SAEN BL77 BL_77 SB77 se_cell
X78 VDD VSS SAEN BL78 BL_78 SB78 se_cell
X79 VDD VSS SAEN BL79 BL_79 SB79 se_cell
X80 VDD VSS SAEN BL80 BL_80 SB80 se_cell
X81 VDD VSS SAEN BL81 BL_81 SB81 se_cell
X82 VDD VSS SAEN BL82 BL_82 SB82 se_cell
X83 VDD VSS SAEN BL83 BL_83 SB83 se_cell
X84 VDD VSS SAEN BL84 BL_84 SB84 se_cell
X85 VDD VSS SAEN BL85 BL_85 SB85 se_cell
X86 VDD VSS SAEN BL86 BL_86 SB86 se_cell
X87 VDD VSS SAEN BL87 BL_87 SB87 se_cell
X88 VDD VSS SAEN BL88 BL_88 SB88 se_cell
X89 VDD VSS SAEN BL89 BL_89 SB89 se_cell
X90 VDD VSS SAEN BL90 BL_90 SB90 se_cell
X91 VDD VSS SAEN BL91 BL_91 SB91 se_cell
X92 VDD VSS SAEN BL92 BL_92 SB92 se_cell
X93 VDD VSS SAEN BL93 BL_93 SB93 se_cell
X94 VDD VSS SAEN BL94 BL_94 SB94 se_cell
X95 VDD VSS SAEN BL95 BL_95 SB95 se_cell
X96 VDD VSS SAEN BL96 BL_96 SB96 se_cell
X97 VDD VSS SAEN BL97 BL_97 SB97 se_cell
X98 VDD VSS SAEN BL98 BL_98 SB98 se_cell
X99 VDD VSS SAEN BL99 BL_99 SB99 se_cell
X100 VDD VSS SAEN BL100 BL_100 SB100 se_cell
X101 VDD VSS SAEN BL101 BL_101 SB101 se_cell
X102 VDD VSS SAEN BL102 BL_102 SB102 se_cell
X103 VDD VSS SAEN BL103 BL_103 SB103 se_cell
X104 VDD VSS SAEN BL104 BL_104 SB104 se_cell
X105 VDD VSS SAEN BL105 BL_105 SB105 se_cell
X106 VDD VSS SAEN BL106 BL_106 SB106 se_cell
X107 VDD VSS SAEN BL107 BL_107 SB107 se_cell
X108 VDD VSS SAEN BL108 BL_108 SB108 se_cell
X109 VDD VSS SAEN BL109 BL_109 SB109 se_cell
X110 VDD VSS SAEN BL110 BL_110 SB110 se_cell
X111 VDD VSS SAEN BL111 BL_111 SB111 se_cell
X112 VDD VSS SAEN BL112 BL_112 SB112 se_cell
X113 VDD VSS SAEN BL113 BL_113 SB113 se_cell
X114 VDD VSS SAEN BL114 BL_114 SB114 se_cell
X115 VDD VSS SAEN BL115 BL_115 SB115 se_cell
X116 VDD VSS SAEN BL116 BL_116 SB116 se_cell
X117 VDD VSS SAEN BL117 BL_117 SB117 se_cell
X118 VDD VSS SAEN BL118 BL_118 SB118 se_cell
X119 VDD VSS SAEN BL119 BL_119 SB119 se_cell
X120 VDD VSS SAEN BL120 BL_120 SB120 se_cell
X121 VDD VSS SAEN BL121 BL_121 SB121 se_cell
X122 VDD VSS SAEN BL122 BL_122 SB122 se_cell
X123 VDD VSS SAEN BL123 BL_123 SB123 se_cell
X124 VDD VSS SAEN BL124 BL_124 SB124 se_cell
X125 VDD VSS SAEN BL125 BL_125 SB125 se_cell
X126 VDD VSS SAEN BL126 BL_126 SB126 se_cell
X127 VDD VSS SAEN BL127 BL_127 SB127 se_cell
.ends se_arr_128

.subckt mat_arr_512 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31
X0 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL0 bit_arr_512
X1 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL1 bit_arr_512
X2 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL2 bit_arr_512
X3 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL3 bit_arr_512
X4 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL4 bit_arr_512
X5 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL5 bit_arr_512
X6 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL6 bit_arr_512
X7 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL7 bit_arr_512
X8 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL8 bit_arr_512
X9 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL9 bit_arr_512
X10 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL10 bit_arr_512
X11 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL11 bit_arr_512
X12 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL12 bit_arr_512
X13 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL13 bit_arr_512
X14 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL14 bit_arr_512
X15 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL15 bit_arr_512
X16 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL16 bit_arr_512
X17 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL17 bit_arr_512
X18 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL18 bit_arr_512
X19 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL19 bit_arr_512
X20 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL20 bit_arr_512
X21 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL21 bit_arr_512
X22 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL22 bit_arr_512
X23 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL23 bit_arr_512
X24 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL24 bit_arr_512
X25 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL25 bit_arr_512
X26 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL26 bit_arr_512
X27 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL27 bit_arr_512
X28 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL28 bit_arr_512
X29 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL29 bit_arr_512
X30 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL30 bit_arr_512
X31 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL31 bit_arr_512
.ends mat_arr_512

.subckt sram128x128 VDD VSS clk addr0 addr1 addr2 addr3 addr4 addr5 addr6 din0 din1 din2 din3 din4 din5 din6 din7 din8 din9 din10 din11 din12 din13 din14 din15 din16 din17 din18 din19 din20 din21 din22 din23 din24 din25 din26 din27 din28 din29 din30 din31 din32 din33 din34 din35 din36 din37 din38 din39 din40 din41 din42 din43 din44 din45 din46 din47 din48 din49 din50 din51 din52 din53 din54 din55 din56 din57 din58 din59 din60 din61 din62 din63 din64 din65 din66 din67 din68 din69 din70 din71 din72 din73 din74 din75 din76 din77 din78 din79 din80 din81 din82 din83 din84 din85 din86 din87 din88 din89 din90 din91 din92 din93 din94 din95 din96 din97 din98 din99 din100 din101 din102 din103 din104 din105 din106 din107 din108 din109 din110 din111 din112 din113 din114 din115 din116 din117 din118 din119 din120 din121 din122 din123 din124 din125 din126 din127 Q0 Q1 Q2 Q3 Q4 Q5 Q6 Q7 Q8 Q9 Q10 Q11 Q12 Q13 Q14 Q15 Q16 Q17 Q18 Q19 Q20 Q21 Q22 Q23 Q24 Q25 Q26 Q27 Q28 Q29 Q30 Q31 Q32 Q33 Q34 Q35 Q36 Q37 Q38 Q39 Q40 Q41 Q42 Q43 Q44 Q45 Q46 Q47 Q48 Q49 Q50 Q51 Q52 Q53 Q54 Q55 Q56 Q57 Q58 Q59 Q60 Q61 Q62 Q63 Q64 Q65 Q66 Q67 Q68 Q69 Q70 Q71 Q72 Q73 Q74 Q75 Q76 Q77 Q78 Q79 Q80 Q81 Q82 Q83 Q84 Q85 Q86 Q87 Q88 Q89 Q90 Q91 Q92 Q93 Q94 Q95 Q96 Q97 Q98 Q99 Q100 Q101 Q102 Q103 Q104 Q105 Q106 Q107 Q108 Q109 Q110 Q111 Q112 Q113 Q114 Q115 Q116 Q117 Q118 Q119 Q120 Q121 Q122 Q123 Q124 Q125 Q126 Q127 w_en cs
X0 VDD VSS clk addr0 addr1 addr2 addr3 addr4 addr5 addr6 w_en A0 A1 A2 A3 A4 A5 A6 write input_reg8
X1 VDD VSS A2 A3 A4 A5 A6 DC0 DC1 DC2 DC3 DC4 DC5 DC6 DC7 DC8 DC9 DC10 DC11 DC12 DC13 DC14 DC15 DC16 DC17 DC18 DC19 DC20 DC21 DC22 DC23 DC24 DC25 DC26 DC27 DC28 DC29 DC30 DC31 row_dec32
X2 VDD VSS WLEN DC0 DC1 DC2 DC3 DC4 DC5 DC6 DC7 DC8 DC9 DC10 DC11 DC12 DC13 DC14 DC15 DC16 DC17 DC18 DC19 DC20 DC21 DC22 DC23 DC24 DC25 DC26 DC27 DC28 DC29 DC30 DC31 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 rd_arr_32
X3 VDD VSS A0 A1 CD0 CD1 CD2 CD3 col_dec4
X4 VDD VSS WLEN CD0 CD1 CD2 CD3 SEL0 SEL1 SEL2 SEL3 rd_arr_4
X5 VDD VSS PCHG WREN SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 SEL0 SEL1 SEL2 SEL3 BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 DW0 DW_0 DW0 DW_0 DW0 DW_0 DW0 DW_0 DW1 DW_1 DW1 DW_1 DW1 DW_1 DW1 DW_1 DW2 DW_2 DW2 DW_2 DW2 DW_2 DW2 DW_2 DW3 DW_3 DW3 DW_3 DW3 DW_3 DW3 DW_3 DW4 DW_4 DW4 DW_4 DW4 DW_4 DW4 DW_4 DW5 DW_5 DW5 DW_5 DW5 DW_5 DW5 DW_5 DW6 DW_6 DW6 DW_6 DW6 DW_6 DW6 DW_6 DW7 DW_7 DW7 DW_7 DW7 DW_7 DW7 DW_7 DW8 DW_8 DW8 DW_8 DW8 DW_8 DW8 DW_8 DW9 DW_9 DW9 DW_9 DW9 DW_9 DW9 DW_9 DW10 DW_10 DW10 DW_10 DW10 DW_10 DW10 DW_10 DW11 DW_11 DW11 DW_11 DW11 DW_11 DW11 DW_11 DW12 DW_12 DW12 DW_12 DW12 DW_12 DW12 DW_12 DW13 DW_13 DW13 DW_13 DW13 DW_13 DW13 DW_13 DW14 DW_14 DW14 DW_14 DW14 DW_14 DW14 DW_14 DW15 DW_15 DW15 DW_15 DW15 DW_15 DW15 DW_15 DW16 DW_16 DW16 DW_16 DW16 DW_16 DW16 DW_16 DW17 DW_17 DW17 DW_17 DW17 DW_17 DW17 DW_17 DW18 DW_18 DW18 DW_18 DW18 DW_18 DW18 DW_18 DW19 DW_19 DW19 DW_19 DW19 DW_19 DW19 DW_19 DW20 DW_20 DW20 DW_20 DW20 DW_20 DW20 DW_20 DW21 DW_21 DW21 DW_21 DW21 DW_21 DW21 DW_21 DW22 DW_22 DW22 DW_22 DW22 DW_22 DW22 DW_22 DW23 DW_23 DW23 DW_23 DW23 DW_23 DW23 DW_23 DW24 DW_24 DW24 DW_24 DW24 DW_24 DW24 DW_24 DW25 DW_25 DW25 DW_25 DW25 DW_25 DW25 DW_25 DW26 DW_26 DW26 DW_26 DW26 DW_26 DW26 DW_26 DW27 DW_27 DW27 DW_27 DW27 DW_27 DW27 DW_27 DW28 DW_28 DW28 DW_28 DW28 DW_28 DW28 DW_28 DW29 DW_29 DW29 DW_29 DW29 DW_29 DW29 DW_29 DW30 DW_30 DW30 DW_30 DW30 DW_30 DW30 DW_30 DW31 DW_31 DW31 DW_31 DW31 DW_31 DW31 DW_31 DW32 DW_32 DW32 DW_32 DW32 DW_32 DW32 DW_32 DW33 DW_33 DW33 DW_33 DW33 DW_33 DW33 DW_33 DW34 DW_34 DW34 DW_34 DW34 DW_34 DW34 DW_34 DW35 DW_35 DW35 DW_35 DW35 DW_35 DW35 DW_35 DW36 DW_36 DW36 DW_36 DW36 DW_36 DW36 DW_36 DW37 DW_37 DW37 DW_37 DW37 DW_37 DW37 DW_37 DW38 DW_38 DW38 DW_38 DW38 DW_38 DW38 DW_38 DW39 DW_39 DW39 DW_39 DW39 DW_39 DW39 DW_39 DW40 DW_40 DW40 DW_40 DW40 DW_40 DW40 DW_40 DW41 DW_41 DW41 DW_41 DW41 DW_41 DW41 DW_41 DW42 DW_42 DW42 DW_42 DW42 DW_42 DW42 DW_42 DW43 DW_43 DW43 DW_43 DW43 DW_43 DW43 DW_43 DW44 DW_44 DW44 DW_44 DW44 DW_44 DW44 DW_44 DW45 DW_45 DW45 DW_45 DW45 DW_45 DW45 DW_45 DW46 DW_46 DW46 DW_46 DW46 DW_46 DW46 DW_46 DW47 DW_47 DW47 DW_47 DW47 DW_47 DW47 DW_47 DW48 DW_48 DW48 DW_48 DW48 DW_48 DW48 DW_48 DW49 DW_49 DW49 DW_49 DW49 DW_49 DW49 DW_49 DW50 DW_50 DW50 DW_50 DW50 DW_50 DW50 DW_50 DW51 DW_51 DW51 DW_51 DW51 DW_51 DW51 DW_51 DW52 DW_52 DW52 DW_52 DW52 DW_52 DW52 DW_52 DW53 DW_53 DW53 DW_53 DW53 DW_53 DW53 DW_53 DW54 DW_54 DW54 DW_54 DW54 DW_54 DW54 DW_54 DW55 DW_55 DW55 DW_55 DW55 DW_55 DW55 DW_55 DW56 DW_56 DW56 DW_56 DW56 DW_56 DW56 DW_56 DW57 DW_57 DW57 DW_57 DW57 DW_57 DW57 DW_57 DW58 DW_58 DW58 DW_58 DW58 DW_58 DW58 DW_58 DW59 DW_59 DW59 DW_59 DW59 DW_59 DW59 DW_59 DW60 DW_60 DW60 DW_60 DW60 DW_60 DW60 DW_60 DW61 DW_61 DW61 DW_61 DW61 DW_61 DW61 DW_61 DW62 DW_62 DW62 DW_62 DW62 DW_62 DW62 DW_62 DW63 DW_63 DW63 DW_63 DW63 DW_63 DW63 DW_63 DW64 DW_64 DW64 DW_64 DW64 DW_64 DW64 DW_64 DW65 DW_65 DW65 DW_65 DW65 DW_65 DW65 DW_65 DW66 DW_66 DW66 DW_66 DW66 DW_66 DW66 DW_66 DW67 DW_67 DW67 DW_67 DW67 DW_67 DW67 DW_67 DW68 DW_68 DW68 DW_68 DW68 DW_68 DW68 DW_68 DW69 DW_69 DW69 DW_69 DW69 DW_69 DW69 DW_69 DW70 DW_70 DW70 DW_70 DW70 DW_70 DW70 DW_70 DW71 DW_71 DW71 DW_71 DW71 DW_71 DW71 DW_71 DW72 DW_72 DW72 DW_72 DW72 DW_72 DW72 DW_72 DW73 DW_73 DW73 DW_73 DW73 DW_73 DW73 DW_73 DW74 DW_74 DW74 DW_74 DW74 DW_74 DW74 DW_74 DW75 DW_75 DW75 DW_75 DW75 DW_75 DW75 DW_75 DW76 DW_76 DW76 DW_76 DW76 DW_76 DW76 DW_76 DW77 DW_77 DW77 DW_77 DW77 DW_77 DW77 DW_77 DW78 DW_78 DW78 DW_78 DW78 DW_78 DW78 DW_78 DW79 DW_79 DW79 DW_79 DW79 DW_79 DW79 DW_79 DW80 DW_80 DW80 DW_80 DW80 DW_80 DW80 DW_80 DW81 DW_81 DW81 DW_81 DW81 DW_81 DW81 DW_81 DW82 DW_82 DW82 DW_82 DW82 DW_82 DW82 DW_82 DW83 DW_83 DW83 DW_83 DW83 DW_83 DW83 DW_83 DW84 DW_84 DW84 DW_84 DW84 DW_84 DW84 DW_84 DW85 DW_85 DW85 DW_85 DW85 DW_85 DW85 DW_85 DW86 DW_86 DW86 DW_86 DW86 DW_86 DW86 DW_86 DW87 DW_87 DW87 DW_87 DW87 DW_87 DW87 DW_87 DW88 DW_88 DW88 DW_88 DW88 DW_88 DW88 DW_88 DW89 DW_89 DW89 DW_89 DW89 DW_89 DW89 DW_89 DW90 DW_90 DW90 DW_90 DW90 DW_90 DW90 DW_90 DW91 DW_91 DW91 DW_91 DW91 DW_91 DW91 DW_91 DW92 DW_92 DW92 DW_92 DW92 DW_92 DW92 DW_92 DW93 DW_93 DW93 DW_93 DW93 DW_93 DW93 DW_93 DW94 DW_94 DW94 DW_94 DW94 DW_94 DW94 DW_94 DW95 DW_95 DW95 DW_95 DW95 DW_95 DW95 DW_95 DW96 DW_96 DW96 DW_96 DW96 DW_96 DW96 DW_96 DW97 DW_97 DW97 DW_97 DW97 DW_97 DW97 DW_97 DW98 DW_98 DW98 DW_98 DW98 DW_98 DW98 DW_98 DW99 DW_99 DW99 DW_99 DW99 DW_99 DW99 DW_99 DW100 DW_100 DW100 DW_100 DW100 DW_100 DW100 DW_100 DW101 DW_101 DW101 DW_101 DW101 DW_101 DW101 DW_101 DW102 DW_102 DW102 DW_102 DW102 DW_102 DW102 DW_102 DW103 DW_103 DW103 DW_103 DW103 DW_103 DW103 DW_103 DW104 DW_104 DW104 DW_104 DW104 DW_104 DW104 DW_104 DW105 DW_105 DW105 DW_105 DW105 DW_105 DW105 DW_105 DW106 DW_106 DW106 DW_106 DW106 DW_106 DW106 DW_106 DW107 DW_107 DW107 DW_107 DW107 DW_107 DW107 DW_107 DW108 DW_108 DW108 DW_108 DW108 DW_108 DW108 DW_108 DW109 DW_109 DW109 DW_109 DW109 DW_109 DW109 DW_109 DW110 DW_110 DW110 DW_110 DW110 DW_110 DW110 DW_110 DW111 DW_111 DW111 DW_111 DW111 DW_111 DW111 DW_111 DW112 DW_112 DW112 DW_112 DW112 DW_112 DW112 DW_112 DW113 DW_113 DW113 DW_113 DW113 DW_113 DW113 DW_113 DW114 DW_114 DW114 DW_114 DW114 DW_114 DW114 DW_114 DW115 DW_115 DW115 DW_115 DW115 DW_115 DW115 DW_115 DW116 DW_116 DW116 DW_116 DW116 DW_116 DW116 DW_116 DW117 DW_117 DW117 DW_117 DW117 DW_117 DW117 DW_117 DW118 DW_118 DW118 DW_118 DW118 DW_118 DW118 DW_118 DW119 DW_119 DW119 DW_119 DW119 DW_119 DW119 DW_119 DW120 DW_120 DW120 DW_120 DW120 DW_120 DW120 DW_120 DW121 DW_121 DW121 DW_121 DW121 DW_121 DW121 DW_121 DW122 DW_122 DW122 DW_122 DW122 DW_122 DW122 DW_122 DW123 DW_123 DW123 DW_123 DW123 DW_123 DW123 DW_123 DW124 DW_124 DW124 DW_124 DW124 DW_124 DW124 DW_124 DW125 DW_125 DW125 DW_125 DW125 DW_125 DW125 DW_125 DW126 DW_126 DW126 DW_126 DW126 DW_126 DW126 DW_126 DW127 DW_127 DW127 DW_127 DW127 DW_127 DW127 DW_127 DR0 DR_0 DR0 DR_0 DR0 DR_0 DR0 DR_0 DR1 DR_1 DR1 DR_1 DR1 DR_1 DR1 DR_1 DR2 DR_2 DR2 DR_2 DR2 DR_2 DR2 DR_2 DR3 DR_3 DR3 DR_3 DR3 DR_3 DR3 DR_3 DR4 DR_4 DR4 DR_4 DR4 DR_4 DR4 DR_4 DR5 DR_5 DR5 DR_5 DR5 DR_5 DR5 DR_5 DR6 DR_6 DR6 DR_6 DR6 DR_6 DR6 DR_6 DR7 DR_7 DR7 DR_7 DR7 DR_7 DR7 DR_7 DR8 DR_8 DR8 DR_8 DR8 DR_8 DR8 DR_8 DR9 DR_9 DR9 DR_9 DR9 DR_9 DR9 DR_9 DR10 DR_10 DR10 DR_10 DR10 DR_10 DR10 DR_10 DR11 DR_11 DR11 DR_11 DR11 DR_11 DR11 DR_11 DR12 DR_12 DR12 DR_12 DR12 DR_12 DR12 DR_12 DR13 DR_13 DR13 DR_13 DR13 DR_13 DR13 DR_13 DR14 DR_14 DR14 DR_14 DR14 DR_14 DR14 DR_14 DR15 DR_15 DR15 DR_15 DR15 DR_15 DR15 DR_15 DR16 DR_16 DR16 DR_16 DR16 DR_16 DR16 DR_16 DR17 DR_17 DR17 DR_17 DR17 DR_17 DR17 DR_17 DR18 DR_18 DR18 DR_18 DR18 DR_18 DR18 DR_18 DR19 DR_19 DR19 DR_19 DR19 DR_19 DR19 DR_19 DR20 DR_20 DR20 DR_20 DR20 DR_20 DR20 DR_20 DR21 DR_21 DR21 DR_21 DR21 DR_21 DR21 DR_21 DR22 DR_22 DR22 DR_22 DR22 DR_22 DR22 DR_22 DR23 DR_23 DR23 DR_23 DR23 DR_23 DR23 DR_23 DR24 DR_24 DR24 DR_24 DR24 DR_24 DR24 DR_24 DR25 DR_25 DR25 DR_25 DR25 DR_25 DR25 DR_25 DR26 DR_26 DR26 DR_26 DR26 DR_26 DR26 DR_26 DR27 DR_27 DR27 DR_27 DR27 DR_27 DR27 DR_27 DR28 DR_28 DR28 DR_28 DR28 DR_28 DR28 DR_28 DR29 DR_29 DR29 DR_29 DR29 DR_29 DR29 DR_29 DR30 DR_30 DR30 DR_30 DR30 DR_30 DR30 DR_30 DR31 DR_31 DR31 DR_31 DR31 DR_31 DR31 DR_31 DR32 DR_32 DR32 DR_32 DR32 DR_32 DR32 DR_32 DR33 DR_33 DR33 DR_33 DR33 DR_33 DR33 DR_33 DR34 DR_34 DR34 DR_34 DR34 DR_34 DR34 DR_34 DR35 DR_35 DR35 DR_35 DR35 DR_35 DR35 DR_35 DR36 DR_36 DR36 DR_36 DR36 DR_36 DR36 DR_36 DR37 DR_37 DR37 DR_37 DR37 DR_37 DR37 DR_37 DR38 DR_38 DR38 DR_38 DR38 DR_38 DR38 DR_38 DR39 DR_39 DR39 DR_39 DR39 DR_39 DR39 DR_39 DR40 DR_40 DR40 DR_40 DR40 DR_40 DR40 DR_40 DR41 DR_41 DR41 DR_41 DR41 DR_41 DR41 DR_41 DR42 DR_42 DR42 DR_42 DR42 DR_42 DR42 DR_42 DR43 DR_43 DR43 DR_43 DR43 DR_43 DR43 DR_43 DR44 DR_44 DR44 DR_44 DR44 DR_44 DR44 DR_44 DR45 DR_45 DR45 DR_45 DR45 DR_45 DR45 DR_45 DR46 DR_46 DR46 DR_46 DR46 DR_46 DR46 DR_46 DR47 DR_47 DR47 DR_47 DR47 DR_47 DR47 DR_47 DR48 DR_48 DR48 DR_48 DR48 DR_48 DR48 DR_48 DR49 DR_49 DR49 DR_49 DR49 DR_49 DR49 DR_49 DR50 DR_50 DR50 DR_50 DR50 DR_50 DR50 DR_50 DR51 DR_51 DR51 DR_51 DR51 DR_51 DR51 DR_51 DR52 DR_52 DR52 DR_52 DR52 DR_52 DR52 DR_52 DR53 DR_53 DR53 DR_53 DR53 DR_53 DR53 DR_53 DR54 DR_54 DR54 DR_54 DR54 DR_54 DR54 DR_54 DR55 DR_55 DR55 DR_55 DR55 DR_55 DR55 DR_55 DR56 DR_56 DR56 DR_56 DR56 DR_56 DR56 DR_56 DR57 DR_57 DR57 DR_57 DR57 DR_57 DR57 DR_57 DR58 DR_58 DR58 DR_58 DR58 DR_58 DR58 DR_58 DR59 DR_59 DR59 DR_59 DR59 DR_59 DR59 DR_59 DR60 DR_60 DR60 DR_60 DR60 DR_60 DR60 DR_60 DR61 DR_61 DR61 DR_61 DR61 DR_61 DR61 DR_61 DR62 DR_62 DR62 DR_62 DR62 DR_62 DR62 DR_62 DR63 DR_63 DR63 DR_63 DR63 DR_63 DR63 DR_63 DR64 DR_64 DR64 DR_64 DR64 DR_64 DR64 DR_64 DR65 DR_65 DR65 DR_65 DR65 DR_65 DR65 DR_65 DR66 DR_66 DR66 DR_66 DR66 DR_66 DR66 DR_66 DR67 DR_67 DR67 DR_67 DR67 DR_67 DR67 DR_67 DR68 DR_68 DR68 DR_68 DR68 DR_68 DR68 DR_68 DR69 DR_69 DR69 DR_69 DR69 DR_69 DR69 DR_69 DR70 DR_70 DR70 DR_70 DR70 DR_70 DR70 DR_70 DR71 DR_71 DR71 DR_71 DR71 DR_71 DR71 DR_71 DR72 DR_72 DR72 DR_72 DR72 DR_72 DR72 DR_72 DR73 DR_73 DR73 DR_73 DR73 DR_73 DR73 DR_73 DR74 DR_74 DR74 DR_74 DR74 DR_74 DR74 DR_74 DR75 DR_75 DR75 DR_75 DR75 DR_75 DR75 DR_75 DR76 DR_76 DR76 DR_76 DR76 DR_76 DR76 DR_76 DR77 DR_77 DR77 DR_77 DR77 DR_77 DR77 DR_77 DR78 DR_78 DR78 DR_78 DR78 DR_78 DR78 DR_78 DR79 DR_79 DR79 DR_79 DR79 DR_79 DR79 DR_79 DR80 DR_80 DR80 DR_80 DR80 DR_80 DR80 DR_80 DR81 DR_81 DR81 DR_81 DR81 DR_81 DR81 DR_81 DR82 DR_82 DR82 DR_82 DR82 DR_82 DR82 DR_82 DR83 DR_83 DR83 DR_83 DR83 DR_83 DR83 DR_83 DR84 DR_84 DR84 DR_84 DR84 DR_84 DR84 DR_84 DR85 DR_85 DR85 DR_85 DR85 DR_85 DR85 DR_85 DR86 DR_86 DR86 DR_86 DR86 DR_86 DR86 DR_86 DR87 DR_87 DR87 DR_87 DR87 DR_87 DR87 DR_87 DR88 DR_88 DR88 DR_88 DR88 DR_88 DR88 DR_88 DR89 DR_89 DR89 DR_89 DR89 DR_89 DR89 DR_89 DR90 DR_90 DR90 DR_90 DR90 DR_90 DR90 DR_90 DR91 DR_91 DR91 DR_91 DR91 DR_91 DR91 DR_91 DR92 DR_92 DR92 DR_92 DR92 DR_92 DR92 DR_92 DR93 DR_93 DR93 DR_93 DR93 DR_93 DR93 DR_93 DR94 DR_94 DR94 DR_94 DR94 DR_94 DR94 DR_94 DR95 DR_95 DR95 DR_95 DR95 DR_95 DR95 DR_95 DR96 DR_96 DR96 DR_96 DR96 DR_96 DR96 DR_96 DR97 DR_97 DR97 DR_97 DR97 DR_97 DR97 DR_97 DR98 DR_98 DR98 DR_98 DR98 DR_98 DR98 DR_98 DR99 DR_99 DR99 DR_99 DR99 DR_99 DR99 DR_99 DR100 DR_100 DR100 DR_100 DR100 DR_100 DR100 DR_100 DR101 DR_101 DR101 DR_101 DR101 DR_101 DR101 DR_101 DR102 DR_102 DR102 DR_102 DR102 DR_102 DR102 DR_102 DR103 DR_103 DR103 DR_103 DR103 DR_103 DR103 DR_103 DR104 DR_104 DR104 DR_104 DR104 DR_104 DR104 DR_104 DR105 DR_105 DR105 DR_105 DR105 DR_105 DR105 DR_105 DR106 DR_106 DR106 DR_106 DR106 DR_106 DR106 DR_106 DR107 DR_107 DR107 DR_107 DR107 DR_107 DR107 DR_107 DR108 DR_108 DR108 DR_108 DR108 DR_108 DR108 DR_108 DR109 DR_109 DR109 DR_109 DR109 DR_109 DR109 DR_109 DR110 DR_110 DR110 DR_110 DR110 DR_110 DR110 DR_110 DR111 DR_111 DR111 DR_111 DR111 DR_111 DR111 DR_111 DR112 DR_112 DR112 DR_112 DR112 DR_112 DR112 DR_112 DR113 DR_113 DR113 DR_113 DR113 DR_113 DR113 DR_113 DR114 DR_114 DR114 DR_114 DR114 DR_114 DR114 DR_114 DR115 DR_115 DR115 DR_115 DR115 DR_115 DR115 DR_115 DR116 DR_116 DR116 DR_116 DR116 DR_116 DR116 DR_116 DR117 DR_117 DR117 DR_117 DR117 DR_117 DR117 DR_117 DR118 DR_118 DR118 DR_118 DR118 DR_118 DR118 DR_118 DR119 DR_119 DR119 DR_119 DR119 DR_119 DR119 DR_119 DR120 DR_120 DR120 DR_120 DR120 DR_120 DR120 DR_120 DR121 DR_121 DR121 DR_121 DR121 DR_121 DR121 DR_121 DR122 DR_122 DR122 DR_122 DR122 DR_122 DR122 DR_122 DR123 DR_123 DR123 DR_123 DR123 DR_123 DR123 DR_123 DR124 DR_124 DR124 DR_124 DR124 DR_124 DR124 DR_124 DR125 DR_125 DR125 DR_125 DR125 DR_125 DR125 DR_125 DR126 DR_126 DR126 DR_126 DR126 DR_126 DR126 DR_126 DR127 DR_127 DR127 DR_127 DR127 DR_127 DR127 DR_127 dido_arr_512
X6 VDD VSS clk WREN din0 din1 din2 din3 din4 din5 din6 din7 din8 din9 din10 din11 din12 din13 din14 din15 din16 din17 din18 din19 din20 din21 din22 din23 din24 din25 din26 din27 din28 din29 din30 din31 din32 din33 din34 din35 din36 din37 din38 din39 din40 din41 din42 din43 din44 din45 din46 din47 din48 din49 din50 din51 din52 din53 din54 din55 din56 din57 din58 din59 din60 din61 din62 din63 din64 din65 din66 din67 din68 din69 din70 din71 din72 din73 din74 din75 din76 din77 din78 din79 din80 din81 din82 din83 din84 din85 din86 din87 din88 din89 din90 din91 din92 din93 din94 din95 din96 din97 din98 din99 din100 din101 din102 din103 din104 din105 din106 din107 din108 din109 din110 din111 din112 din113 din114 din115 din116 din117 din118 din119 din120 din121 din122 din123 din124 din125 din126 din127 DW0 DW_0 DW1 DW_1 DW2 DW_2 DW3 DW_3 DW4 DW_4 DW5 DW_5 DW6 DW_6 DW7 DW_7 DW8 DW_8 DW9 DW_9 DW10 DW_10 DW11 DW_11 DW12 DW_12 DW13 DW_13 DW14 DW_14 DW15 DW_15 DW16 DW_16 DW17 DW_17 DW18 DW_18 DW19 DW_19 DW20 DW_20 DW21 DW_21 DW22 DW_22 DW23 DW_23 DW24 DW_24 DW25 DW_25 DW26 DW_26 DW27 DW_27 DW28 DW_28 DW29 DW_29 DW30 DW_30 DW31 DW_31 DW32 DW_32 DW33 DW_33 DW34 DW_34 DW35 DW_35 DW36 DW_36 DW37 DW_37 DW38 DW_38 DW39 DW_39 DW40 DW_40 DW41 DW_41 DW42 DW_42 DW43 DW_43 DW44 DW_44 DW45 DW_45 DW46 DW_46 DW47 DW_47 DW48 DW_48 DW49 DW_49 DW50 DW_50 DW51 DW_51 DW52 DW_52 DW53 DW_53 DW54 DW_54 DW55 DW_55 DW56 DW_56 DW57 DW_57 DW58 DW_58 DW59 DW_59 DW60 DW_60 DW61 DW_61 DW62 DW_62 DW63 DW_63 DW64 DW_64 DW65 DW_65 DW66 DW_66 DW67 DW_67 DW68 DW_68 DW69 DW_69 DW70 DW_70 DW71 DW_71 DW72 DW_72 DW73 DW_73 DW74 DW_74 DW75 DW_75 DW76 DW_76 DW77 DW_77 DW78 DW_78 DW79 DW_79 DW80 DW_80 DW81 DW_81 DW82 DW_82 DW83 DW_83 DW84 DW_84 DW85 DW_85 DW86 DW_86 DW87 DW_87 DW88 DW_88 DW89 DW_89 DW90 DW_90 DW91 DW_91 DW92 DW_92 DW93 DW_93 DW94 DW_94 DW95 DW_95 DW96 DW_96 DW97 DW_97 DW98 DW_98 DW99 DW_99 DW100 DW_100 DW101 DW_101 DW102 DW_102 DW103 DW_103 DW104 DW_104 DW105 DW_105 DW106 DW_106 DW107 DW_107 DW108 DW_108 DW109 DW_109 DW110 DW_110 DW111 DW_111 DW112 DW_112 DW113 DW_113 DW114 DW_114 DW115 DW_115 DW116 DW_116 DW117 DW_117 DW118 DW_118 DW119 DW_119 DW120 DW_120 DW121 DW_121 DW122 DW_122 DW123 DW_123 DW124 DW_124 DW125 DW_125 DW126 DW_126 DW127 DW_127 datain_reg128
X7 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 BL64 BL_64 BL65 BL_65 BL66 BL_66 BL67 BL_67 BL68 BL_68 BL69 BL_69 BL70 BL_70 BL71 BL_71 BL72 BL_72 BL73 BL_73 BL74 BL_74 BL75 BL_75 BL76 BL_76 BL77 BL_77 BL78 BL_78 BL79 BL_79 BL80 BL_80 BL81 BL_81 BL82 BL_82 BL83 BL_83 BL84 BL_84 BL85 BL_85 BL86 BL_86 BL87 BL_87 BL88 BL_88 BL89 BL_89 BL90 BL_90 BL91 BL_91 BL92 BL_92 BL93 BL_93 BL94 BL_94 BL95 BL_95 BL96 BL_96 BL97 BL_97 BL98 BL_98 BL99 BL_99 BL100 BL_100 BL101 BL_101 BL102 BL_102 BL103 BL_103 BL104 BL_104 BL105 BL_105 BL106 BL_106 BL107 BL_107 BL108 BL_108 BL109 BL_109 BL110 BL_110 BL111 BL_111 BL112 BL_112 BL113 BL_113 BL114 BL_114 BL115 BL_115 BL116 BL_116 BL117 BL_117 BL118 BL_118 BL119 BL_119 BL120 BL_120 BL121 BL_121 BL122 BL_122 BL123 BL_123 BL124 BL_124 BL125 BL_125 BL126 BL_126 BL127 BL_127 BL128 BL_128 BL129 BL_129 BL130 BL_130 BL131 BL_131 BL132 BL_132 BL133 BL_133 BL134 BL_134 BL135 BL_135 BL136 BL_136 BL137 BL_137 BL138 BL_138 BL139 BL_139 BL140 BL_140 BL141 BL_141 BL142 BL_142 BL143 BL_143 BL144 BL_144 BL145 BL_145 BL146 BL_146 BL147 BL_147 BL148 BL_148 BL149 BL_149 BL150 BL_150 BL151 BL_151 BL152 BL_152 BL153 BL_153 BL154 BL_154 BL155 BL_155 BL156 BL_156 BL157 BL_157 BL158 BL_158 BL159 BL_159 BL160 BL_160 BL161 BL_161 BL162 BL_162 BL163 BL_163 BL164 BL_164 BL165 BL_165 BL166 BL_166 BL167 BL_167 BL168 BL_168 BL169 BL_169 BL170 BL_170 BL171 BL_171 BL172 BL_172 BL173 BL_173 BL174 BL_174 BL175 BL_175 BL176 BL_176 BL177 BL_177 BL178 BL_178 BL179 BL_179 BL180 BL_180 BL181 BL_181 BL182 BL_182 BL183 BL_183 BL184 BL_184 BL185 BL_185 BL186 BL_186 BL187 BL_187 BL188 BL_188 BL189 BL_189 BL190 BL_190 BL191 BL_191 BL192 BL_192 BL193 BL_193 BL194 BL_194 BL195 BL_195 BL196 BL_196 BL197 BL_197 BL198 BL_198 BL199 BL_199 BL200 BL_200 BL201 BL_201 BL202 BL_202 BL203 BL_203 BL204 BL_204 BL205 BL_205 BL206 BL_206 BL207 BL_207 BL208 BL_208 BL209 BL_209 BL210 BL_210 BL211 BL_211 BL212 BL_212 BL213 BL_213 BL214 BL_214 BL215 BL_215 BL216 BL_216 BL217 BL_217 BL218 BL_218 BL219 BL_219 BL220 BL_220 BL221 BL_221 BL222 BL_222 BL223 BL_223 BL224 BL_224 BL225 BL_225 BL226 BL_226 BL227 BL_227 BL228 BL_228 BL229 BL_229 BL230 BL_230 BL231 BL_231 BL232 BL_232 BL233 BL_233 BL234 BL_234 BL235 BL_235 BL236 BL_236 BL237 BL_237 BL238 BL_238 BL239 BL_239 BL240 BL_240 BL241 BL_241 BL242 BL_242 BL243 BL_243 BL244 BL_244 BL245 BL_245 BL246 BL_246 BL247 BL_247 BL248 BL_248 BL249 BL_249 BL250 BL_250 BL251 BL_251 BL252 BL_252 BL253 BL_253 BL254 BL_254 BL255 BL_255 BL256 BL_256 BL257 BL_257 BL258 BL_258 BL259 BL_259 BL260 BL_260 BL261 BL_261 BL262 BL_262 BL263 BL_263 BL264 BL_264 BL265 BL_265 BL266 BL_266 BL267 BL_267 BL268 BL_268 BL269 BL_269 BL270 BL_270 BL271 BL_271 BL272 BL_272 BL273 BL_273 BL274 BL_274 BL275 BL_275 BL276 BL_276 BL277 BL_277 BL278 BL_278 BL279 BL_279 BL280 BL_280 BL281 BL_281 BL282 BL_282 BL283 BL_283 BL284 BL_284 BL285 BL_285 BL286 BL_286 BL287 BL_287 BL288 BL_288 BL289 BL_289 BL290 BL_290 BL291 BL_291 BL292 BL_292 BL293 BL_293 BL294 BL_294 BL295 BL_295 BL296 BL_296 BL297 BL_297 BL298 BL_298 BL299 BL_299 BL300 BL_300 BL301 BL_301 BL302 BL_302 BL303 BL_303 BL304 BL_304 BL305 BL_305 BL306 BL_306 BL307 BL_307 BL308 BL_308 BL309 BL_309 BL310 BL_310 BL311 BL_311 BL312 BL_312 BL313 BL_313 BL314 BL_314 BL315 BL_315 BL316 BL_316 BL317 BL_317 BL318 BL_318 BL319 BL_319 BL320 BL_320 BL321 BL_321 BL322 BL_322 BL323 BL_323 BL324 BL_324 BL325 BL_325 BL326 BL_326 BL327 BL_327 BL328 BL_328 BL329 BL_329 BL330 BL_330 BL331 BL_331 BL332 BL_332 BL333 BL_333 BL334 BL_334 BL335 BL_335 BL336 BL_336 BL337 BL_337 BL338 BL_338 BL339 BL_339 BL340 BL_340 BL341 BL_341 BL342 BL_342 BL343 BL_343 BL344 BL_344 BL345 BL_345 BL346 BL_346 BL347 BL_347 BL348 BL_348 BL349 BL_349 BL350 BL_350 BL351 BL_351 BL352 BL_352 BL353 BL_353 BL354 BL_354 BL355 BL_355 BL356 BL_356 BL357 BL_357 BL358 BL_358 BL359 BL_359 BL360 BL_360 BL361 BL_361 BL362 BL_362 BL363 BL_363 BL364 BL_364 BL365 BL_365 BL366 BL_366 BL367 BL_367 BL368 BL_368 BL369 BL_369 BL370 BL_370 BL371 BL_371 BL372 BL_372 BL373 BL_373 BL374 BL_374 BL375 BL_375 BL376 BL_376 BL377 BL_377 BL378 BL_378 BL379 BL_379 BL380 BL_380 BL381 BL_381 BL382 BL_382 BL383 BL_383 BL384 BL_384 BL385 BL_385 BL386 BL_386 BL387 BL_387 BL388 BL_388 BL389 BL_389 BL390 BL_390 BL391 BL_391 BL392 BL_392 BL393 BL_393 BL394 BL_394 BL395 BL_395 BL396 BL_396 BL397 BL_397 BL398 BL_398 BL399 BL_399 BL400 BL_400 BL401 BL_401 BL402 BL_402 BL403 BL_403 BL404 BL_404 BL405 BL_405 BL406 BL_406 BL407 BL_407 BL408 BL_408 BL409 BL_409 BL410 BL_410 BL411 BL_411 BL412 BL_412 BL413 BL_413 BL414 BL_414 BL415 BL_415 BL416 BL_416 BL417 BL_417 BL418 BL_418 BL419 BL_419 BL420 BL_420 BL421 BL_421 BL422 BL_422 BL423 BL_423 BL424 BL_424 BL425 BL_425 BL426 BL_426 BL427 BL_427 BL428 BL_428 BL429 BL_429 BL430 BL_430 BL431 BL_431 BL432 BL_432 BL433 BL_433 BL434 BL_434 BL435 BL_435 BL436 BL_436 BL437 BL_437 BL438 BL_438 BL439 BL_439 BL440 BL_440 BL441 BL_441 BL442 BL_442 BL443 BL_443 BL444 BL_444 BL445 BL_445 BL446 BL_446 BL447 BL_447 BL448 BL_448 BL449 BL_449 BL450 BL_450 BL451 BL_451 BL452 BL_452 BL453 BL_453 BL454 BL_454 BL455 BL_455 BL456 BL_456 BL457 BL_457 BL458 BL_458 BL459 BL_459 BL460 BL_460 BL461 BL_461 BL462 BL_462 BL463 BL_463 BL464 BL_464 BL465 BL_465 BL466 BL_466 BL467 BL_467 BL468 BL_468 BL469 BL_469 BL470 BL_470 BL471 BL_471 BL472 BL_472 BL473 BL_473 BL474 BL_474 BL475 BL_475 BL476 BL_476 BL477 BL_477 BL478 BL_478 BL479 BL_479 BL480 BL_480 BL481 BL_481 BL482 BL_482 BL483 BL_483 BL484 BL_484 BL485 BL_485 BL486 BL_486 BL487 BL_487 BL488 BL_488 BL489 BL_489 BL490 BL_490 BL491 BL_491 BL492 BL_492 BL493 BL_493 BL494 BL_494 BL495 BL_495 BL496 BL_496 BL497 BL_497 BL498 BL_498 BL499 BL_499 BL500 BL_500 BL501 BL_501 BL502 BL_502 BL503 BL_503 BL504 BL_504 BL505 BL_505 BL506 BL_506 BL507 BL_507 BL508 BL_508 BL509 BL_509 BL510 BL_510 BL511 BL_511 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 mat_arr_512
X8 VDD VSS SAEN DR0 DR_0 DR1 DR_1 DR2 DR_2 DR3 DR_3 DR4 DR_4 DR5 DR_5 DR6 DR_6 DR7 DR_7 DR8 DR_8 DR9 DR_9 DR10 DR_10 DR11 DR_11 DR12 DR_12 DR13 DR_13 DR14 DR_14 DR15 DR_15 DR16 DR_16 DR17 DR_17 DR18 DR_18 DR19 DR_19 DR20 DR_20 DR21 DR_21 DR22 DR_22 DR23 DR_23 DR24 DR_24 DR25 DR_25 DR26 DR_26 DR27 DR_27 DR28 DR_28 DR29 DR_29 DR30 DR_30 DR31 DR_31 DR32 DR_32 DR33 DR_33 DR34 DR_34 DR35 DR_35 DR36 DR_36 DR37 DR_37 DR38 DR_38 DR39 DR_39 DR40 DR_40 DR41 DR_41 DR42 DR_42 DR43 DR_43 DR44 DR_44 DR45 DR_45 DR46 DR_46 DR47 DR_47 DR48 DR_48 DR49 DR_49 DR50 DR_50 DR51 DR_51 DR52 DR_52 DR53 DR_53 DR54 DR_54 DR55 DR_55 DR56 DR_56 DR57 DR_57 DR58 DR_58 DR59 DR_59 DR60 DR_60 DR61 DR_61 DR62 DR_62 DR63 DR_63 DR64 DR_64 DR65 DR_65 DR66 DR_66 DR67 DR_67 DR68 DR_68 DR69 DR_69 DR70 DR_70 DR71 DR_71 DR72 DR_72 DR73 DR_73 DR74 DR_74 DR75 DR_75 DR76 DR_76 DR77 DR_77 DR78 DR_78 DR79 DR_79 DR80 DR_80 DR81 DR_81 DR82 DR_82 DR83 DR_83 DR84 DR_84 DR85 DR_85 DR86 DR_86 DR87 DR_87 DR88 DR_88 DR89 DR_89 DR90 DR_90 DR91 DR_91 DR92 DR_92 DR93 DR_93 DR94 DR_94 DR95 DR_95 DR96 DR_96 DR97 DR_97 DR98 DR_98 DR99 DR_99 DR100 DR_100 DR101 DR_101 DR102 DR_102 DR103 DR_103 DR104 DR_104 DR105 DR_105 DR106 DR_106 DR107 DR_107 DR108 DR_108 DR109 DR_109 DR110 DR_110 DR111 DR_111 DR112 DR_112 DR113 DR_113 DR114 DR_114 DR115 DR_115 DR116 DR_116 DR117 DR_117 DR118 DR_118 DR119 DR_119 DR120 DR_120 DR121 DR_121 DR122 DR_122 DR123 DR_123 DR124 DR_124 DR125 DR_125 DR126 DR_126 DR127 DR_127 Q0 Q1 Q2 Q3 Q4 Q5 Q6 Q7 Q8 Q9 Q10 Q11 Q12 Q13 Q14 Q15 Q16 Q17 Q18 Q19 Q20 Q21 Q22 Q23 Q24 Q25 Q26 Q27 Q28 Q29 Q30 Q31 Q32 Q33 Q34 Q35 Q36 Q37 Q38 Q39 Q40 Q41 Q42 Q43 Q44 Q45 Q46 Q47 Q48 Q49 Q50 Q51 Q52 Q53 Q54 Q55 Q56 Q57 Q58 Q59 Q60 Q61 Q62 Q63 Q64 Q65 Q66 Q67 Q68 Q69 Q70 Q71 Q72 Q73 Q74 Q75 Q76 Q77 Q78 Q79 Q80 Q81 Q82 Q83 Q84 Q85 Q86 Q87 Q88 Q89 Q90 Q91 Q92 Q93 Q94 Q95 Q96 Q97 Q98 Q99 Q100 Q101 Q102 Q103 Q104 Q105 Q106 Q107 Q108 Q109 Q110 Q111 Q112 Q113 Q114 Q115 Q116 Q117 Q118 Q119 Q120 Q121 Q122 Q123 Q124 Q125 Q126 Q127 se_arr_128
X9 VDD VSS clk cs write DBL DBL_ WREN PCHG WLEN SAEN ctrl
X10 VDD VSS WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 DBL DBL_ dmy_arr_32
.ends sram128x128

