magic
tech sky130A
magscale 1 2
timestamp 1703576186
<< nwell >>
rect 1711 1541 3864 1749
rect 2820 1144 3038 1541
rect 3395 1540 3864 1541
rect 3428 1144 3864 1540
rect 1711 936 3864 1144
rect 3088 935 3864 936
rect 3176 825 3864 935
rect 3176 620 3394 825
<< pwell >>
rect 1721 1364 1831 1376
rect 2433 1364 2543 1376
rect 1721 1228 2031 1364
rect 2433 1228 2743 1364
rect 1721 1216 1831 1228
rect 2433 1216 2543 1228
rect 3076 1364 3186 1376
rect 3076 1228 3386 1364
rect 3076 1216 3186 1228
rect 2462 759 2572 771
rect 2462 623 2772 759
rect 2462 611 2572 623
<< nmos >>
rect 1917 1254 1947 1338
rect 2211 1254 2241 1338
rect 2299 1254 2329 1338
rect 2629 1254 2659 1338
rect 3272 1254 3302 1338
rect 1805 648 1835 732
rect 2023 648 2053 732
rect 2240 649 2270 733
rect 2328 649 2358 733
rect 2658 649 2688 733
rect 2876 649 2906 733
rect 2964 649 2994 733
rect 3270 349 3300 549
rect 3522 349 3552 749
rect 3740 349 3770 749
<< pmos >>
rect 1917 1603 1947 1687
rect 2211 1603 2241 1687
rect 2299 1603 2329 1687
rect 2629 1603 2659 1687
rect 2870 1603 2900 1687
rect 2958 1603 2988 1687
rect 3272 1603 3302 1687
rect 2914 1389 2944 1473
rect 1805 998 1835 1082
rect 2023 998 2053 1082
rect 2240 998 2270 1082
rect 2328 998 2358 1082
rect 2658 998 2688 1082
rect 2876 998 2906 1082
rect 2964 998 2994 1082
rect 3270 682 3300 1082
rect 3522 887 3552 1687
rect 3740 887 3770 1687
<< ndiff >>
rect 1859 1313 1917 1338
rect 1859 1279 1871 1313
rect 1905 1279 1917 1313
rect 1859 1254 1917 1279
rect 1947 1313 2005 1338
rect 1947 1279 1959 1313
rect 1993 1279 2005 1313
rect 1947 1254 2005 1279
rect 2153 1326 2211 1338
rect 2153 1266 2165 1326
rect 2199 1266 2211 1326
rect 2153 1254 2211 1266
rect 2241 1326 2299 1338
rect 2241 1266 2253 1326
rect 2287 1266 2299 1326
rect 2241 1254 2299 1266
rect 2329 1326 2387 1338
rect 2329 1266 2341 1326
rect 2375 1266 2387 1326
rect 2329 1254 2387 1266
rect 2571 1313 2629 1338
rect 2571 1279 2583 1313
rect 2617 1279 2629 1313
rect 2571 1254 2629 1279
rect 2659 1313 2717 1338
rect 2659 1279 2671 1313
rect 2705 1279 2717 1313
rect 2659 1254 2717 1279
rect 3214 1313 3272 1338
rect 3214 1279 3226 1313
rect 3260 1279 3272 1313
rect 3214 1254 3272 1279
rect 3302 1313 3360 1338
rect 3302 1279 3314 1313
rect 3348 1279 3360 1313
rect 3302 1254 3360 1279
rect 1747 720 1805 732
rect 1747 660 1759 720
rect 1793 660 1805 720
rect 1747 648 1805 660
rect 1835 720 1893 732
rect 1835 660 1847 720
rect 1881 660 1893 720
rect 1835 648 1893 660
rect 1965 720 2023 732
rect 1965 660 1977 720
rect 2011 660 2023 720
rect 1965 648 2023 660
rect 2053 720 2111 732
rect 2053 660 2065 720
rect 2099 660 2111 720
rect 2053 648 2111 660
rect 2182 721 2240 733
rect 2182 661 2194 721
rect 2228 661 2240 721
rect 2182 649 2240 661
rect 2270 721 2328 733
rect 2270 661 2282 721
rect 2316 661 2328 721
rect 2270 649 2328 661
rect 2358 721 2416 733
rect 2358 661 2370 721
rect 2404 661 2416 721
rect 2358 649 2416 661
rect 2600 708 2658 733
rect 2600 674 2612 708
rect 2646 674 2658 708
rect 2600 649 2658 674
rect 2688 708 2746 733
rect 2688 674 2700 708
rect 2734 674 2746 708
rect 2688 649 2746 674
rect 2818 721 2876 733
rect 2818 661 2830 721
rect 2864 661 2876 721
rect 2818 649 2876 661
rect 2906 721 2964 733
rect 2906 661 2918 721
rect 2952 661 2964 721
rect 2906 649 2964 661
rect 2994 721 3052 733
rect 2994 661 3006 721
rect 3040 661 3052 721
rect 3464 737 3522 749
rect 2994 649 3052 661
rect 3212 537 3270 549
rect 3212 361 3224 537
rect 3258 361 3270 537
rect 3212 349 3270 361
rect 3300 537 3358 549
rect 3300 361 3312 537
rect 3346 361 3358 537
rect 3300 349 3358 361
rect 3464 361 3476 737
rect 3510 361 3522 737
rect 3464 349 3522 361
rect 3552 737 3610 749
rect 3552 361 3564 737
rect 3598 361 3610 737
rect 3552 349 3610 361
rect 3682 737 3740 749
rect 3682 361 3694 737
rect 3728 361 3740 737
rect 3682 349 3740 361
rect 3770 737 3828 749
rect 3770 361 3782 737
rect 3816 361 3828 737
rect 3770 349 3828 361
<< pdiff >>
rect 1859 1662 1917 1687
rect 1859 1628 1871 1662
rect 1905 1628 1917 1662
rect 1859 1603 1917 1628
rect 1947 1662 2005 1687
rect 1947 1628 1959 1662
rect 1993 1628 2005 1662
rect 1947 1603 2005 1628
rect 2153 1675 2211 1687
rect 2153 1615 2165 1675
rect 2199 1615 2211 1675
rect 2153 1603 2211 1615
rect 2241 1675 2299 1687
rect 2241 1615 2253 1675
rect 2287 1615 2299 1675
rect 2241 1603 2299 1615
rect 2329 1675 2387 1687
rect 2329 1615 2341 1675
rect 2375 1615 2387 1675
rect 2329 1603 2387 1615
rect 2571 1662 2629 1687
rect 2571 1628 2583 1662
rect 2617 1628 2629 1662
rect 2571 1603 2629 1628
rect 2659 1662 2717 1687
rect 2659 1628 2671 1662
rect 2705 1628 2717 1662
rect 2659 1603 2717 1628
rect 2812 1675 2870 1687
rect 2812 1615 2824 1675
rect 2858 1615 2870 1675
rect 2812 1603 2870 1615
rect 2900 1675 2958 1687
rect 2900 1615 2912 1675
rect 2946 1615 2958 1675
rect 2900 1603 2958 1615
rect 2988 1675 3046 1687
rect 2988 1615 3000 1675
rect 3034 1615 3046 1675
rect 2988 1603 3046 1615
rect 3214 1662 3272 1687
rect 3214 1628 3226 1662
rect 3260 1628 3272 1662
rect 3214 1603 3272 1628
rect 3302 1662 3360 1687
rect 3302 1628 3314 1662
rect 3348 1628 3360 1662
rect 3302 1603 3360 1628
rect 3464 1675 3522 1687
rect 2856 1461 2914 1473
rect 2856 1401 2868 1461
rect 2902 1401 2914 1461
rect 2856 1389 2914 1401
rect 2944 1461 3002 1473
rect 2944 1401 2956 1461
rect 2990 1401 3002 1461
rect 2944 1389 3002 1401
rect 1747 1070 1805 1082
rect 1747 1010 1759 1070
rect 1793 1010 1805 1070
rect 1747 998 1805 1010
rect 1835 1070 1893 1082
rect 1835 1010 1847 1070
rect 1881 1010 1893 1070
rect 1835 998 1893 1010
rect 1965 1070 2023 1082
rect 1965 1010 1977 1070
rect 2011 1010 2023 1070
rect 1965 998 2023 1010
rect 2053 1070 2111 1082
rect 2053 1010 2065 1070
rect 2099 1010 2111 1070
rect 2053 998 2111 1010
rect 2182 1070 2240 1082
rect 2182 1010 2194 1070
rect 2228 1010 2240 1070
rect 2182 998 2240 1010
rect 2270 1070 2328 1082
rect 2270 1010 2282 1070
rect 2316 1010 2328 1070
rect 2270 998 2328 1010
rect 2358 1070 2416 1082
rect 2358 1010 2370 1070
rect 2404 1010 2416 1070
rect 2358 998 2416 1010
rect 2600 1057 2658 1082
rect 2600 1023 2612 1057
rect 2646 1023 2658 1057
rect 2600 998 2658 1023
rect 2688 1057 2746 1082
rect 2688 1023 2700 1057
rect 2734 1023 2746 1057
rect 2688 998 2746 1023
rect 2818 1070 2876 1082
rect 2818 1010 2830 1070
rect 2864 1010 2876 1070
rect 2818 998 2876 1010
rect 2906 1070 2964 1082
rect 2906 1010 2918 1070
rect 2952 1010 2964 1070
rect 2906 998 2964 1010
rect 2994 1070 3052 1082
rect 2994 1010 3006 1070
rect 3040 1010 3052 1070
rect 2994 998 3052 1010
rect 3212 1070 3270 1082
rect 3212 694 3224 1070
rect 3258 694 3270 1070
rect 3212 682 3270 694
rect 3300 1070 3358 1082
rect 3300 694 3312 1070
rect 3346 694 3358 1070
rect 3464 899 3476 1675
rect 3510 899 3522 1675
rect 3464 887 3522 899
rect 3552 1675 3610 1687
rect 3552 899 3564 1675
rect 3598 899 3610 1675
rect 3552 887 3610 899
rect 3682 1675 3740 1687
rect 3682 899 3694 1675
rect 3728 899 3740 1675
rect 3682 887 3740 899
rect 3770 1675 3828 1687
rect 3770 899 3782 1675
rect 3816 899 3828 1675
rect 3770 887 3828 899
rect 3300 682 3358 694
<< ndiffc >>
rect 1871 1279 1905 1313
rect 1959 1279 1993 1313
rect 2165 1266 2199 1326
rect 2253 1266 2287 1326
rect 2341 1266 2375 1326
rect 2583 1279 2617 1313
rect 2671 1279 2705 1313
rect 3226 1279 3260 1313
rect 3314 1279 3348 1313
rect 1759 660 1793 720
rect 1847 660 1881 720
rect 1977 660 2011 720
rect 2065 660 2099 720
rect 2194 661 2228 721
rect 2282 661 2316 721
rect 2370 661 2404 721
rect 2612 674 2646 708
rect 2700 674 2734 708
rect 2830 661 2864 721
rect 2918 661 2952 721
rect 3006 661 3040 721
rect 3224 361 3258 537
rect 3312 361 3346 537
rect 3476 361 3510 737
rect 3564 361 3598 737
rect 3694 361 3728 737
rect 3782 361 3816 737
<< pdiffc >>
rect 1871 1628 1905 1662
rect 1959 1628 1993 1662
rect 2165 1615 2199 1675
rect 2253 1615 2287 1675
rect 2341 1615 2375 1675
rect 2583 1628 2617 1662
rect 2671 1628 2705 1662
rect 2824 1615 2858 1675
rect 2912 1615 2946 1675
rect 3000 1615 3034 1675
rect 3226 1628 3260 1662
rect 3314 1628 3348 1662
rect 2868 1401 2902 1461
rect 2956 1401 2990 1461
rect 1759 1010 1793 1070
rect 1847 1010 1881 1070
rect 1977 1010 2011 1070
rect 2065 1010 2099 1070
rect 2194 1010 2228 1070
rect 2282 1010 2316 1070
rect 2370 1010 2404 1070
rect 2612 1023 2646 1057
rect 2700 1023 2734 1057
rect 2830 1010 2864 1070
rect 2918 1010 2952 1070
rect 3006 1010 3040 1070
rect 3224 694 3258 1070
rect 3312 694 3346 1070
rect 3476 899 3510 1675
rect 3564 899 3598 1675
rect 3694 899 3728 1675
rect 3782 899 3816 1675
<< psubdiff >>
rect 1747 1313 1805 1350
rect 1747 1279 1759 1313
rect 1793 1279 1805 1313
rect 1747 1242 1805 1279
rect 2459 1313 2517 1350
rect 2459 1279 2471 1313
rect 2505 1279 2517 1313
rect 2459 1242 2517 1279
rect 3102 1313 3160 1350
rect 3102 1279 3114 1313
rect 3148 1279 3160 1313
rect 3102 1242 3160 1279
rect 2488 708 2546 745
rect 2488 674 2500 708
rect 2534 674 2546 708
rect 2488 637 2546 674
<< nsubdiff >>
rect 1747 1662 1805 1699
rect 1747 1628 1759 1662
rect 1793 1628 1805 1662
rect 1747 1591 1805 1628
rect 2459 1662 2517 1699
rect 2459 1628 2471 1662
rect 2505 1628 2517 1662
rect 2459 1591 2517 1628
rect 3102 1662 3160 1699
rect 3102 1628 3114 1662
rect 3148 1628 3160 1662
rect 3102 1591 3160 1628
rect 2488 1057 2546 1094
rect 2488 1023 2500 1057
rect 2534 1023 2546 1057
rect 2488 986 2546 1023
<< psubdiffcont >>
rect 1759 1279 1793 1313
rect 2471 1279 2505 1313
rect 3114 1279 3148 1313
rect 2500 674 2534 708
<< nsubdiffcont >>
rect 1759 1628 1793 1662
rect 2471 1628 2505 1662
rect 3114 1628 3148 1662
rect 2500 1023 2534 1057
<< poly >>
rect 1917 1687 1947 1713
rect 2211 1687 2241 1713
rect 2299 1687 2329 1713
rect 2629 1687 2659 1713
rect 2870 1687 2900 1713
rect 2958 1687 2988 1713
rect 1917 1513 1947 1603
rect 2211 1571 2241 1603
rect 1856 1497 1947 1513
rect 2161 1555 2241 1571
rect 2161 1521 2177 1555
rect 2211 1521 2241 1555
rect 2161 1505 2241 1521
rect 1856 1463 1872 1497
rect 1906 1463 1947 1497
rect 1856 1447 1947 1463
rect 1917 1338 1947 1447
rect 2211 1338 2241 1505
rect 2299 1426 2329 1603
rect 3272 1687 3302 1713
rect 3522 1687 3552 1713
rect 3740 1687 3770 1713
rect 2629 1513 2659 1603
rect 2870 1577 2900 1603
rect 2958 1577 2988 1603
rect 2870 1555 2988 1577
rect 2870 1547 2912 1555
rect 2568 1497 2659 1513
rect 2896 1521 2912 1547
rect 2946 1547 2988 1555
rect 2946 1521 2961 1547
rect 2896 1505 2961 1521
rect 3272 1513 3302 1603
rect 2913 1499 2944 1505
rect 2568 1463 2584 1497
rect 2618 1463 2659 1497
rect 2914 1473 2944 1499
rect 3211 1497 3302 1513
rect 2568 1447 2659 1463
rect 2299 1410 2379 1426
rect 2299 1376 2329 1410
rect 2363 1376 2379 1410
rect 2299 1360 2379 1376
rect 2299 1338 2329 1360
rect 2629 1338 2659 1447
rect 3211 1463 3227 1497
rect 3261 1463 3302 1497
rect 3211 1447 3302 1463
rect 2914 1363 2944 1389
rect 1917 1228 1947 1254
rect 2211 1228 2241 1254
rect 2299 1228 2329 1254
rect 3272 1338 3302 1447
rect 2629 1228 2659 1254
rect 3272 1228 3302 1254
rect 1805 1082 1835 1108
rect 2023 1082 2053 1108
rect 2240 1082 2270 1108
rect 2328 1082 2358 1108
rect 2658 1082 2688 1108
rect 2876 1082 2906 1108
rect 2964 1082 2994 1108
rect 3270 1082 3300 1108
rect 1805 935 1835 998
rect 1734 918 1835 935
rect 1734 884 1751 918
rect 1785 884 1835 918
rect 1734 868 1835 884
rect 1805 732 1835 868
rect 2023 832 2053 998
rect 2240 966 2270 998
rect 2190 950 2270 966
rect 2190 916 2206 950
rect 2240 916 2270 950
rect 2190 900 2270 916
rect 1951 816 2053 832
rect 1951 782 1967 816
rect 2001 782 2053 816
rect 1951 766 2053 782
rect 2023 732 2053 766
rect 2240 733 2270 900
rect 2328 821 2358 998
rect 2658 908 2688 998
rect 2876 966 2906 998
rect 2597 892 2688 908
rect 2826 950 2906 966
rect 2826 916 2842 950
rect 2876 916 2906 950
rect 2826 900 2906 916
rect 2597 858 2613 892
rect 2647 858 2688 892
rect 2597 842 2688 858
rect 2328 805 2408 821
rect 2328 771 2358 805
rect 2392 771 2408 805
rect 2328 755 2408 771
rect 2328 733 2358 755
rect 2658 733 2688 842
rect 2876 733 2906 900
rect 2964 821 2994 998
rect 2964 805 3044 821
rect 2964 771 2994 805
rect 3028 771 3044 805
rect 2964 755 3044 771
rect 2964 733 2994 755
rect 1805 622 1835 648
rect 2023 622 2053 648
rect 2240 623 2270 649
rect 2328 623 2358 649
rect 3522 854 3552 887
rect 3740 855 3770 887
rect 3460 838 3552 854
rect 3460 804 3476 838
rect 3510 804 3552 838
rect 3460 788 3552 804
rect 3681 839 3770 855
rect 3681 805 3698 839
rect 3732 805 3770 839
rect 3681 789 3770 805
rect 3522 749 3552 788
rect 3740 749 3770 789
rect 2658 623 2688 649
rect 2876 623 2906 649
rect 2964 623 2994 649
rect 3270 644 3300 682
rect 3208 628 3300 644
rect 3208 594 3224 628
rect 3258 594 3300 628
rect 3208 578 3300 594
rect 3270 549 3300 578
rect 3270 323 3300 349
rect 3522 323 3552 349
rect 3740 323 3770 349
<< polycont >>
rect 2177 1521 2211 1555
rect 1872 1463 1906 1497
rect 2912 1521 2946 1555
rect 2584 1463 2618 1497
rect 2329 1376 2363 1410
rect 3227 1463 3261 1497
rect 1751 884 1785 918
rect 2206 916 2240 950
rect 1967 782 2001 816
rect 2842 916 2876 950
rect 2613 858 2647 892
rect 2358 771 2392 805
rect 2994 771 3028 805
rect 3476 804 3510 838
rect 3698 805 3732 839
rect 3224 594 3258 628
<< locali >>
rect 1747 1662 1905 1691
rect 1747 1628 1759 1662
rect 1793 1628 1871 1662
rect 1747 1599 1905 1628
rect 1959 1662 1993 1691
rect 1959 1497 1993 1628
rect 2165 1675 2199 1691
rect 2165 1599 2199 1615
rect 2253 1675 2287 1691
rect 2253 1599 2287 1615
rect 2341 1675 2375 1691
rect 2341 1599 2375 1615
rect 2459 1662 2617 1691
rect 2459 1628 2471 1662
rect 2505 1628 2583 1662
rect 2459 1599 2617 1628
rect 2671 1662 2705 1691
rect 2161 1521 2177 1555
rect 2211 1521 2227 1555
rect 2671 1497 2705 1628
rect 1856 1463 1872 1497
rect 1906 1463 1922 1497
rect 2568 1463 2584 1497
rect 2618 1463 2634 1497
rect 1759 1313 1905 1342
rect 1793 1279 1871 1313
rect 1759 1250 1905 1279
rect 1959 1313 1993 1463
rect 1959 1250 1993 1279
rect 2063 1376 2177 1410
rect 2211 1376 2329 1410
rect 2363 1376 2379 1410
rect 2063 1178 2097 1376
rect 2165 1326 2199 1342
rect 2165 1250 2199 1266
rect 2253 1326 2287 1342
rect 2253 1250 2287 1266
rect 2341 1326 2375 1342
rect 2341 1250 2375 1266
rect 2471 1313 2617 1342
rect 2505 1279 2583 1313
rect 2471 1250 2617 1279
rect 2671 1313 2705 1463
rect 2824 1675 2858 1691
rect 2824 1483 2858 1615
rect 2912 1675 2946 1691
rect 2912 1599 2946 1615
rect 3000 1675 3034 1691
rect 3000 1599 3034 1615
rect 3102 1662 3260 1691
rect 3102 1628 3114 1662
rect 3148 1628 3226 1662
rect 3102 1599 3260 1628
rect 3314 1662 3348 1691
rect 2896 1521 2912 1555
rect 2946 1521 3130 1555
rect 2824 1461 2902 1483
rect 2824 1449 2868 1461
rect 2868 1385 2902 1401
rect 2956 1461 2990 1477
rect 2956 1385 2990 1401
rect 3096 1429 3130 1521
rect 3314 1497 3348 1628
rect 3211 1463 3227 1497
rect 3261 1463 3277 1497
rect 2671 1250 2705 1279
rect 3114 1313 3260 1342
rect 3148 1279 3226 1313
rect 3114 1250 3260 1279
rect 3314 1313 3348 1463
rect 1847 1144 2097 1178
rect 3314 1170 3348 1279
rect 1759 1070 1793 1086
rect 1759 994 1793 1010
rect 1847 1070 1881 1144
rect 3114 1136 3348 1170
rect 3476 1675 3510 1691
rect 1734 884 1751 918
rect 1785 884 1801 918
rect 1847 816 1881 1010
rect 1977 1070 2011 1086
rect 1977 994 2011 1010
rect 2065 1070 2099 1086
rect 2065 950 2099 1010
rect 2194 1070 2228 1086
rect 2194 994 2228 1010
rect 2282 1070 2316 1086
rect 2282 994 2316 1010
rect 2370 1070 2404 1086
rect 2370 994 2404 1010
rect 2488 1057 2646 1086
rect 2488 1023 2500 1057
rect 2534 1023 2612 1057
rect 2488 994 2646 1023
rect 2700 1057 2734 1086
rect 2065 916 2206 950
rect 2240 916 2256 950
rect 1847 782 1967 816
rect 2001 782 2017 816
rect 1759 720 1793 736
rect 1759 644 1793 660
rect 1847 720 1881 782
rect 1847 644 1881 660
rect 1977 720 2011 736
rect 1977 644 2011 660
rect 2065 720 2099 916
rect 2700 892 2734 1023
rect 2830 1070 2864 1086
rect 2830 994 2864 1010
rect 2918 1070 2952 1086
rect 2918 994 2952 1010
rect 3006 1070 3040 1086
rect 3006 994 3040 1010
rect 2826 916 2842 950
rect 2876 916 2892 950
rect 2597 858 2613 892
rect 2647 858 2663 892
rect 2194 771 2206 805
rect 2240 771 2358 805
rect 2392 771 2408 805
rect 2065 644 2099 660
rect 2194 721 2228 737
rect 2194 645 2228 661
rect 2282 721 2316 737
rect 2282 645 2316 661
rect 2370 721 2404 737
rect 2370 645 2404 661
rect 2500 708 2646 737
rect 2534 674 2612 708
rect 2500 645 2646 674
rect 2700 708 2734 858
rect 3114 805 3148 1136
rect 2830 771 2842 805
rect 2876 771 2994 805
rect 3028 771 3148 805
rect 3224 1070 3258 1086
rect 2700 645 2734 674
rect 2830 721 2864 737
rect 2830 645 2864 661
rect 2918 721 2952 737
rect 2918 645 2952 661
rect 3006 721 3040 737
rect 3224 678 3258 694
rect 3312 1070 3346 1086
rect 3476 883 3510 899
rect 3564 1675 3598 1691
rect 3439 804 3476 838
rect 3510 804 3526 838
rect 3006 628 3040 661
rect 3006 594 3224 628
rect 3258 594 3274 628
rect 3224 537 3258 553
rect 3224 345 3258 361
rect 3312 537 3346 694
rect 3312 345 3346 361
rect 3476 737 3510 753
rect 3476 345 3510 361
rect 3564 737 3598 899
rect 3694 1675 3728 1691
rect 3694 883 3728 899
rect 3782 1675 3816 1691
rect 3687 805 3698 839
rect 3732 805 3748 839
rect 3564 345 3598 361
rect 3694 737 3728 753
rect 3694 345 3728 361
rect 3782 737 3816 899
rect 3782 345 3816 361
<< viali >>
rect 1871 1628 1905 1662
rect 1959 1628 1993 1662
rect 2165 1615 2199 1675
rect 2253 1615 2287 1675
rect 2341 1615 2375 1675
rect 2583 1628 2617 1662
rect 2671 1628 2705 1662
rect 2177 1521 2211 1555
rect 1872 1463 1906 1497
rect 1959 1463 1993 1497
rect 2584 1463 2618 1497
rect 2671 1463 2705 1497
rect 1871 1279 1905 1313
rect 1959 1279 1993 1313
rect 2177 1376 2211 1410
rect 2165 1266 2199 1326
rect 2253 1266 2287 1326
rect 2341 1266 2375 1326
rect 2583 1279 2617 1313
rect 2824 1615 2858 1675
rect 2912 1615 2946 1675
rect 3000 1615 3034 1675
rect 3226 1628 3260 1662
rect 3314 1628 3348 1662
rect 2868 1401 2902 1461
rect 2956 1401 2990 1461
rect 3227 1463 3261 1497
rect 3314 1463 3348 1497
rect 3096 1395 3130 1429
rect 2671 1279 2705 1313
rect 3226 1279 3260 1313
rect 3314 1279 3348 1313
rect 1759 1010 1793 1070
rect 1847 1010 1881 1070
rect 1751 884 1785 918
rect 1977 1010 2011 1070
rect 2065 1010 2099 1070
rect 2194 1010 2228 1070
rect 2282 1010 2316 1070
rect 2370 1010 2404 1070
rect 2612 1023 2646 1057
rect 2700 1023 2734 1057
rect 2206 916 2240 950
rect 1759 660 1793 720
rect 1847 660 1881 720
rect 1977 660 2011 720
rect 2830 1010 2864 1070
rect 2918 1010 2952 1070
rect 3006 1010 3040 1070
rect 2842 916 2876 950
rect 2613 858 2647 892
rect 2700 858 2734 892
rect 2206 771 2240 805
rect 2065 660 2099 720
rect 2194 661 2228 721
rect 2282 661 2316 721
rect 2370 661 2404 721
rect 2612 674 2646 708
rect 2842 771 2876 805
rect 2700 674 2734 708
rect 2830 661 2864 721
rect 2918 661 2952 721
rect 3006 661 3040 721
rect 3224 694 3258 1070
rect 3312 694 3346 1070
rect 3476 899 3510 1675
rect 3564 899 3598 1675
rect 3405 804 3439 838
rect 3224 361 3258 537
rect 3312 361 3346 537
rect 3476 361 3510 737
rect 3694 899 3728 1675
rect 3782 899 3816 1675
rect 3653 805 3687 839
rect 3564 361 3598 737
rect 3694 361 3728 737
rect 3782 361 3816 737
<< metal1 >>
rect 0 1715 3864 1749
rect 1871 1687 1905 1715
rect 2165 1687 2199 1715
rect 2341 1687 2375 1715
rect 2583 1687 2617 1715
rect 2912 1687 2946 1715
rect 3226 1687 3260 1715
rect 3476 1687 3510 1715
rect 3694 1687 3728 1715
rect 1865 1662 1911 1687
rect 1865 1628 1871 1662
rect 1905 1628 1911 1662
rect 1865 1603 1911 1628
rect 1953 1662 1999 1687
rect 1953 1628 1959 1662
rect 1993 1628 1999 1662
rect 1953 1603 1999 1628
rect 2159 1675 2205 1687
rect 2159 1615 2165 1675
rect 2199 1615 2205 1675
rect 2159 1603 2205 1615
rect 2247 1675 2293 1687
rect 2247 1615 2253 1675
rect 2287 1615 2293 1675
rect 2247 1603 2293 1615
rect 2335 1675 2381 1687
rect 2335 1615 2341 1675
rect 2375 1615 2381 1675
rect 2335 1603 2381 1615
rect 2577 1662 2623 1687
rect 2577 1628 2583 1662
rect 2617 1628 2623 1662
rect 2577 1603 2623 1628
rect 2665 1662 2711 1687
rect 2818 1675 2864 1687
rect 2818 1667 2824 1675
rect 2665 1628 2671 1662
rect 2705 1628 2711 1662
rect 2665 1603 2711 1628
rect 2766 1615 2776 1667
rect 2858 1615 2864 1675
rect 2818 1603 2864 1615
rect 2906 1675 2952 1687
rect 2906 1615 2912 1675
rect 2946 1615 2952 1675
rect 2906 1603 2952 1615
rect 2994 1675 3040 1687
rect 2994 1615 3000 1675
rect 3034 1615 3040 1675
rect 3093 1615 3103 1667
rect 3220 1662 3266 1687
rect 3220 1628 3226 1662
rect 3260 1628 3266 1662
rect 2994 1603 3040 1615
rect 3220 1603 3266 1628
rect 3308 1662 3354 1687
rect 3308 1628 3314 1662
rect 3348 1628 3354 1662
rect 3308 1603 3354 1628
rect 3470 1675 3516 1687
rect 2059 1555 2069 1573
rect 2013 1521 2069 1555
rect 2121 1555 2131 1573
rect 2165 1555 2223 1561
rect 2121 1521 2177 1555
rect 2211 1521 2223 1555
rect 2013 1503 2041 1521
rect 2165 1515 2223 1521
rect 1860 1497 1918 1503
rect 0 1463 1872 1497
rect 1906 1463 1918 1497
rect 1860 1457 1918 1463
rect 1947 1497 2041 1503
rect 1947 1463 1959 1497
rect 1993 1463 2041 1497
rect 2253 1497 2287 1603
rect 2572 1497 2630 1503
rect 2253 1463 2584 1497
rect 2618 1463 2630 1497
rect 1947 1457 2005 1463
rect 2165 1410 2223 1416
rect 2117 1376 2177 1410
rect 2211 1376 2223 1410
rect 2165 1370 2223 1376
rect 2341 1338 2375 1463
rect 2572 1457 2630 1463
rect 2659 1497 2717 1503
rect 3000 1497 3034 1603
rect 3215 1497 3273 1503
rect 2659 1463 2671 1497
rect 2705 1463 2787 1497
rect 3000 1473 3227 1497
rect 2659 1457 2717 1463
rect 1865 1313 1911 1338
rect 1865 1279 1871 1313
rect 1905 1279 1911 1313
rect 1865 1254 1911 1279
rect 1953 1313 1999 1338
rect 1953 1279 1959 1313
rect 1993 1279 1999 1313
rect 1953 1254 1999 1279
rect 2159 1326 2205 1338
rect 2159 1266 2165 1326
rect 2199 1266 2205 1326
rect 2159 1254 2205 1266
rect 2247 1326 2293 1338
rect 2247 1266 2253 1326
rect 2287 1266 2293 1326
rect 2247 1254 2293 1266
rect 2335 1326 2381 1338
rect 2335 1266 2341 1326
rect 2375 1266 2381 1326
rect 2335 1254 2381 1266
rect 2577 1313 2623 1338
rect 2577 1279 2583 1313
rect 2617 1279 2623 1313
rect 2577 1254 2623 1279
rect 2665 1313 2711 1338
rect 2665 1279 2671 1313
rect 2705 1279 2711 1313
rect 2753 1301 2787 1463
rect 2862 1461 2908 1473
rect 2862 1401 2868 1461
rect 2902 1401 2908 1461
rect 2862 1389 2908 1401
rect 2950 1463 3227 1473
rect 3261 1463 3273 1497
rect 2950 1461 3034 1463
rect 2950 1401 2956 1461
rect 2990 1435 3034 1461
rect 3215 1457 3273 1463
rect 3302 1497 3360 1503
rect 3302 1463 3314 1497
rect 3348 1463 3396 1497
rect 3302 1457 3360 1463
rect 2990 1401 2996 1435
rect 2950 1389 2996 1401
rect 3084 1429 3142 1435
rect 3084 1395 3096 1429
rect 3130 1425 3142 1429
rect 3130 1395 3376 1425
rect 3084 1389 3376 1395
rect 3366 1373 3376 1389
rect 3428 1373 3438 1425
rect 2839 1301 2849 1353
rect 3220 1313 3266 1338
rect 2665 1254 2711 1279
rect 3220 1279 3226 1313
rect 3260 1279 3266 1313
rect 3220 1254 3266 1279
rect 3308 1313 3354 1338
rect 3308 1279 3314 1313
rect 3348 1279 3354 1313
rect 3308 1254 3354 1279
rect 1871 1225 1905 1254
rect 2165 1225 2199 1254
rect 2583 1225 2617 1254
rect 3226 1225 3260 1254
rect 0 1191 3396 1225
rect 3470 1144 3476 1675
rect 0 1110 3476 1144
rect 1759 1082 1793 1110
rect 1977 1082 2011 1110
rect 2194 1082 2228 1110
rect 2370 1082 2404 1110
rect 2612 1082 2646 1110
rect 2830 1082 2864 1110
rect 3006 1082 3040 1110
rect 3224 1082 3258 1110
rect 1753 1070 1799 1082
rect 1753 1010 1759 1070
rect 1793 1010 1799 1070
rect 1753 998 1799 1010
rect 1841 1070 1887 1082
rect 1841 1010 1847 1070
rect 1881 1010 1887 1070
rect 1841 998 1887 1010
rect 1971 1070 2017 1082
rect 1971 1010 1977 1070
rect 2011 1010 2017 1070
rect 1971 998 2017 1010
rect 2059 1070 2105 1082
rect 2059 1010 2065 1070
rect 2099 1010 2105 1070
rect 2059 998 2105 1010
rect 2188 1070 2234 1082
rect 2188 1010 2194 1070
rect 2228 1010 2234 1070
rect 2188 998 2234 1010
rect 2276 1070 2322 1082
rect 2276 1010 2282 1070
rect 2316 1010 2322 1070
rect 2276 998 2322 1010
rect 2364 1070 2410 1082
rect 2364 1010 2370 1070
rect 2404 1010 2410 1070
rect 2364 998 2410 1010
rect 2606 1057 2652 1082
rect 2606 1023 2612 1057
rect 2646 1023 2652 1057
rect 2606 998 2652 1023
rect 2694 1057 2740 1082
rect 2694 1023 2700 1057
rect 2734 1023 2740 1057
rect 2694 998 2740 1023
rect 2824 1070 2870 1082
rect 2824 1010 2830 1070
rect 2864 1010 2870 1070
rect 2824 998 2870 1010
rect 2912 1070 2958 1082
rect 2912 1010 2918 1070
rect 2952 1010 2958 1070
rect 2912 998 2958 1010
rect 3000 1070 3046 1082
rect 3000 1010 3006 1070
rect 3040 1010 3046 1070
rect 3000 998 3046 1010
rect 3218 1070 3264 1082
rect 2194 950 2252 956
rect 0 891 1522 925
rect 1488 805 1522 891
rect 1602 884 1612 936
rect 1664 918 1674 936
rect 1739 918 1797 924
rect 1664 884 1751 918
rect 1785 884 1797 918
rect 2146 916 2206 950
rect 2240 916 2252 950
rect 2194 910 2252 916
rect 1739 878 1797 884
rect 2282 892 2316 998
rect 2830 950 2888 956
rect 2782 949 2842 950
rect 2748 916 2842 949
rect 2876 916 2888 950
rect 2748 910 2888 916
rect 2748 904 2830 910
rect 2737 898 2747 904
rect 2601 892 2659 898
rect 2282 858 2613 892
rect 2647 858 2659 892
rect 2194 805 2252 811
rect 1488 771 2206 805
rect 2240 771 2252 805
rect 2194 765 2252 771
rect 2370 733 2404 858
rect 2601 852 2659 858
rect 2688 892 2747 898
rect 2688 858 2700 892
rect 2734 858 2747 892
rect 2688 852 2747 858
rect 2799 852 2809 904
rect 2918 892 2952 998
rect 2918 858 3088 892
rect 2830 805 2888 811
rect 2782 771 2842 805
rect 2876 771 2888 805
rect 2830 765 2888 771
rect 3006 733 3040 858
rect 1753 720 1799 732
rect 1753 660 1759 720
rect 1793 660 1799 720
rect 1753 648 1799 660
rect 1841 720 1887 732
rect 1841 660 1847 720
rect 1881 660 1887 720
rect 1841 648 1887 660
rect 1971 720 2017 732
rect 1971 660 1977 720
rect 2011 660 2017 720
rect 1971 648 2017 660
rect 2059 720 2105 732
rect 2059 660 2065 720
rect 2099 660 2105 720
rect 2059 648 2105 660
rect 2188 721 2234 733
rect 2188 661 2194 721
rect 2228 661 2234 721
rect 2188 649 2234 661
rect 2276 721 2322 733
rect 2276 661 2282 721
rect 2316 661 2322 721
rect 2276 649 2322 661
rect 2364 721 2410 733
rect 2364 661 2370 721
rect 2404 661 2410 721
rect 2364 649 2410 661
rect 2606 708 2652 733
rect 2606 674 2612 708
rect 2646 674 2652 708
rect 2606 649 2652 674
rect 2694 708 2740 733
rect 2694 674 2700 708
rect 2734 674 2740 708
rect 2694 649 2740 674
rect 2824 721 2870 733
rect 2824 661 2830 721
rect 2864 661 2870 721
rect 2824 649 2870 661
rect 2912 721 2958 733
rect 2912 661 2918 721
rect 2952 661 2958 721
rect 2912 649 2958 661
rect 3000 721 3046 733
rect 3000 661 3006 721
rect 3040 661 3046 721
rect 3218 694 3224 1070
rect 3258 694 3264 1070
rect 3218 682 3264 694
rect 3306 1070 3352 1082
rect 3306 694 3312 1070
rect 3346 694 3352 1070
rect 3470 899 3476 1110
rect 3510 899 3516 1675
rect 3470 887 3516 899
rect 3558 1675 3604 1687
rect 3558 899 3564 1675
rect 3598 899 3604 1675
rect 3558 887 3604 899
rect 3688 1675 3734 1687
rect 3688 899 3694 1675
rect 3728 899 3734 1675
rect 3688 887 3734 899
rect 3776 1675 3822 1687
rect 3776 899 3782 1675
rect 3816 899 3822 1675
rect 3776 887 3822 899
rect 3388 798 3398 850
rect 3450 798 3460 850
rect 3502 795 3512 847
rect 3564 749 3598 887
rect 3634 798 3644 850
rect 3696 798 3706 850
rect 3782 749 3816 887
rect 4018 759 4316 768
rect 3306 682 3352 694
rect 3470 737 3516 749
rect 3000 649 3046 661
rect 1759 620 1793 648
rect 1977 620 2011 648
rect 2194 620 2228 649
rect 2612 620 2646 649
rect 2830 620 2864 649
rect 0 619 3088 620
rect 0 586 3122 619
rect 1602 503 1612 521
rect 0 469 1612 503
rect 1664 469 1674 521
rect 3088 318 3122 586
rect 3218 537 3264 549
rect 3218 361 3224 537
rect 3258 361 3264 537
rect 3218 349 3264 361
rect 3306 537 3352 549
rect 3306 361 3312 537
rect 3346 361 3352 537
rect 3306 349 3352 361
rect 3470 361 3476 737
rect 3510 361 3516 737
rect 3470 349 3516 361
rect 3558 737 3604 749
rect 3558 361 3564 737
rect 3598 361 3604 737
rect 3558 349 3604 361
rect 3688 737 3734 749
rect 3688 361 3694 737
rect 3728 361 3734 737
rect 3688 349 3734 361
rect 3776 737 3822 749
rect 3776 361 3782 737
rect 3816 361 3822 737
rect 4018 707 4028 759
rect 4081 734 4316 759
rect 4081 707 4091 734
rect 3776 349 3822 361
rect 3224 318 3258 349
rect 3476 318 3510 349
rect 3694 318 3728 349
rect 3088 284 3728 318
rect 3782 34 3816 349
rect 3782 0 4316 34
<< via1 >>
rect 2776 1615 2824 1667
rect 2824 1615 2829 1667
rect 3040 1615 3093 1667
rect 2069 1521 2121 1573
rect 3376 1373 3428 1425
rect 2787 1301 2839 1353
rect 1612 884 1664 936
rect 2747 852 2799 904
rect 3398 838 3450 850
rect 3398 804 3405 838
rect 3405 804 3439 838
rect 3439 804 3450 838
rect 3398 798 3450 804
rect 3512 795 3564 847
rect 3644 839 3696 850
rect 3644 805 3653 839
rect 3653 805 3687 839
rect 3687 805 3696 839
rect 3644 798 3696 805
rect 1612 469 1664 521
rect 4028 707 4081 759
<< metal2 >>
rect 2765 2027 2817 2133
rect 2658 1993 2817 2027
rect 2658 1832 2692 1993
rect 3634 1909 3686 2133
rect 1795 1798 2692 1832
rect 2795 1875 3686 1909
rect 2795 1801 2830 1875
rect 4224 1835 4276 2133
rect 3059 1801 4276 1835
rect 1612 936 1664 946
rect 1612 521 1664 884
rect 1795 876 1829 1798
rect 2795 1677 2829 1801
rect 3059 1677 3093 1801
rect 2776 1667 2829 1677
rect 2776 1605 2829 1615
rect 3040 1667 3093 1677
rect 3040 1605 3093 1615
rect 2069 1573 2121 1583
rect 2069 1512 2121 1521
rect 2069 1477 3644 1512
rect 3376 1425 3428 1435
rect 3428 1373 3546 1406
rect 3376 1363 3546 1373
rect 2787 1353 2839 1363
rect 2839 1301 3398 1325
rect 2787 1291 3398 1301
rect 2747 904 2799 914
rect 1795 852 2747 876
rect 1795 842 2799 852
rect 3364 860 3398 1291
rect 3364 850 3450 860
rect 3364 798 3398 850
rect 3364 788 3450 798
rect 3512 857 3546 1363
rect 3610 860 3644 1477
rect 3512 847 3564 857
rect 3512 785 3564 795
rect 3610 850 3696 860
rect 3610 798 3644 850
rect 3610 788 3696 798
rect 3512 741 3546 785
rect 4028 759 4081 769
rect 3512 707 4028 741
rect 4028 697 4081 707
rect 1612 459 1664 469
<< labels >>
rlabel metal2 2765 2081 2817 2133 0 WLEN
rlabel metal2 3634 2081 3686 2133 0 DBL
rlabel metal2 4224 2081 4276 2133 0 DBL_
rlabel metal1 4282 734 4316 768 0 PCHG
rlabel metal1 4282 0 4316 34 0 WREN
rlabel metal1 0 1715 34 1749 0 VDD
rlabel metal1 0 1463 34 1497 0 write
rlabel metal1 0 1191 34 1225 0 VSS
rlabel metal1 0 1110 34 1144 0 VDD
rlabel metal1 0 891 34 925 0 cs
rlabel metal1 0 586 34 620 0 VSS
rlabel metal1 0 469 34 503 0 clk
<< end >>
