magic
tech sky130A
magscale 1 2
timestamp 1702552054
<< nwell >>
rect -109 -146 109 146
<< pmos >>
rect -15 -84 15 84
<< pdiff >>
rect -73 72 -15 84
rect -73 -72 -61 72
rect -27 -72 -15 72
rect -73 -84 -15 -72
rect 15 72 73 84
rect 15 -72 27 72
rect 61 -72 73 72
rect 15 -84 73 -72
<< pdiffc >>
rect -61 -72 -27 72
rect 27 -72 61 72
<< poly >>
rect -15 84 15 110
rect -15 -110 15 -84
<< locali >>
rect -61 72 -27 88
rect -61 -88 -27 -72
rect 27 72 61 88
rect 27 -88 61 -72
<< viali >>
rect -61 -72 -27 72
rect 27 -72 61 72
<< metal1 >>
rect -67 72 -21 84
rect -67 -72 -61 72
rect -27 -72 -21 72
rect -67 -84 -21 -72
rect 21 72 67 84
rect 21 -72 27 72
rect 61 -72 67 72
rect 21 -84 67 -72
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.84 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
