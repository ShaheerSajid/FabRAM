magic
tech sky130A
magscale 1 2
timestamp 1702458901
<< nwell >>
rect 330 1560 709 1768
rect 330 950 709 1158
<< metal1 >>
rect 637 2302 647 2354
rect 699 2302 709 2354
rect 477 2126 487 2178
rect 539 2160 549 2178
rect 539 2126 711 2160
rect 1299 2059 1309 2111
rect 1361 2059 1371 2111
rect 397 1981 407 2033
rect 459 2015 469 2033
rect 459 1981 709 2015
rect 557 1796 567 1848
rect 619 1830 629 1848
rect 619 1796 709 1830
rect 328 1734 647 1768
rect 637 1716 647 1734
rect 699 1716 709 1768
rect 477 1540 487 1592
rect 539 1574 549 1592
rect 539 1540 709 1574
rect 477 1516 505 1540
rect 1299 1522 1309 1525
rect 0 1482 34 1516
rect 330 1482 505 1516
rect 161 1439 195 1482
rect 1297 1476 1309 1522
rect 1299 1473 1309 1476
rect 1361 1473 1371 1525
rect 477 1439 487 1448
rect 161 1405 487 1439
rect 477 1396 487 1405
rect 539 1396 549 1448
rect 647 1395 709 1429
rect 317 1310 327 1362
rect 379 1344 389 1362
rect 647 1344 681 1395
rect 379 1310 681 1344
rect 557 1244 567 1272
rect 327 1220 567 1244
rect 619 1244 629 1272
rect 619 1220 709 1244
rect 327 1210 709 1220
rect 327 1209 455 1210
rect 257 1124 647 1158
rect 637 1106 647 1124
rect 699 1106 709 1158
rect 477 930 487 982
rect 539 964 549 982
rect 539 930 709 964
rect 1299 912 1309 915
rect 0 872 34 906
rect 257 872 431 906
rect 161 811 195 872
rect 397 837 431 872
rect 1297 866 1309 912
rect 1299 863 1309 866
rect 1361 863 1371 915
rect 161 777 351 811
rect 397 785 407 837
rect 459 819 469 837
rect 459 785 709 819
rect 317 734 351 777
rect 317 682 327 734
rect 379 682 389 734
rect 557 634 567 662
rect 257 610 567 634
rect 619 634 629 662
rect 619 610 709 634
rect 257 600 709 610
rect 637 516 647 568
rect 699 516 709 568
rect 477 340 487 392
rect 539 374 549 392
rect 539 340 709 374
rect 1299 322 1309 325
rect 1297 276 1309 322
rect 1299 273 1309 276
rect 1361 273 1371 325
rect 316 195 326 247
rect 378 229 388 247
rect 378 195 709 229
rect 557 10 567 62
rect 619 44 629 62
rect 619 10 709 44
<< via1 >>
rect 647 2302 699 2354
rect 487 2126 539 2178
rect 1309 2059 1361 2111
rect 407 1981 459 2033
rect 567 1796 619 1848
rect 647 1716 699 1768
rect 487 1540 539 1592
rect 1309 1473 1361 1525
rect 487 1396 539 1448
rect 327 1310 379 1362
rect 567 1220 619 1272
rect 647 1106 699 1158
rect 487 930 539 982
rect 1309 863 1361 915
rect 407 785 459 837
rect 327 682 379 734
rect 567 610 619 662
rect 647 516 699 568
rect 487 340 539 392
rect 1309 273 1361 325
rect 326 195 378 247
rect 567 10 619 62
<< metal2 >>
rect 487 2178 539 2188
rect 407 2033 459 2043
rect 327 1362 379 1372
rect 327 734 379 1310
rect 407 837 459 1981
rect 487 1592 539 2126
rect 487 1534 539 1540
rect 567 1848 619 2422
rect 407 777 459 785
rect 487 1448 539 1456
rect 487 982 539 1396
rect 327 257 379 682
rect 487 392 539 930
rect 487 331 539 340
rect 567 1272 619 1796
rect 567 662 619 1220
rect 326 247 379 257
rect 378 195 379 247
rect 326 185 379 195
rect 567 62 619 610
rect 567 0 619 10
rect 647 2354 699 2422
rect 647 1768 699 2302
rect 1307 2113 1363 2123
rect 1307 2047 1363 2057
rect 647 1158 699 1716
rect 1307 1527 1363 1537
rect 1307 1461 1363 1471
rect 647 568 699 1106
rect 1307 917 1363 927
rect 1307 851 1363 861
rect 647 0 699 516
rect 1307 327 1363 337
rect 1307 261 1363 271
<< via2 >>
rect 1307 2111 1363 2113
rect 1307 2059 1309 2111
rect 1309 2059 1361 2111
rect 1361 2059 1363 2111
rect 1307 2057 1363 2059
rect 1307 1525 1363 1527
rect 1307 1473 1309 1525
rect 1309 1473 1361 1525
rect 1361 1473 1363 1525
rect 1307 1471 1363 1473
rect 1307 915 1363 917
rect 1307 863 1309 915
rect 1309 863 1361 915
rect 1361 863 1363 915
rect 1307 861 1363 863
rect 1307 325 1363 327
rect 1307 273 1309 325
rect 1309 273 1361 325
rect 1361 273 1363 325
rect 1307 271 1363 273
<< metal3 >>
rect 1297 2113 1462 2118
rect 1297 2057 1307 2113
rect 1363 2057 1462 2113
rect 1297 2052 1462 2057
rect 1297 1527 1462 1532
rect 1297 1471 1307 1527
rect 1363 1471 1462 1527
rect 1297 1466 1462 1471
rect 1297 917 1462 922
rect 1297 861 1307 917
rect 1363 861 1462 917
rect 1297 856 1462 861
rect 1297 327 1462 332
rect 1297 271 1307 327
rect 1363 271 1462 327
rect 1297 266 1462 271
use nand2  nand2_0 ~/Desktop/FabRAM/FE/sram130/nand2
timestamp 1702458901
transform 1 0 709 0 1 1705
box 0 91 306 649
use nand2  nand2_1
timestamp 1702458901
transform 1 0 709 0 1 1119
box 0 91 306 649
use nand2  nand2_2
timestamp 1702458901
transform 1 0 709 0 1 509
box 0 91 306 649
use nand2  nand2_3
timestamp 1702458901
transform 1 0 709 0 1 -81
box 0 91 306 649
use not  not_0 ~/Desktop/FabRAM/FE/sram130/not
timestamp 1702458901
transform 1 0 1015 0 1 1705
box 0 91 330 649
use not  not_1
timestamp 1702458901
transform 1 0 1015 0 1 1119
box 0 91 330 649
use not  not_2
timestamp 1702458901
transform 1 0 1015 0 1 509
box 0 91 330 649
use not  not_3
timestamp 1702458901
transform 1 0 1015 0 1 -81
box 0 91 330 649
use not  not_5
timestamp 1702458901
transform 1 0 0 0 1 509
box 0 91 330 649
use not  not_6
timestamp 1702458901
transform 1 0 0 0 1 1119
box 0 91 330 649
<< labels >>
rlabel metal3 1396 2052 1462 2118 0 Y0
rlabel metal3 1396 1466 1462 1532 0 Y1
rlabel metal3 1396 856 1462 922 0 Y2
rlabel metal3 1396 266 1462 332 0 Y3
rlabel metal2 567 2370 619 2422 0 VSS
rlabel metal2 647 2370 699 2422 0 VDD
rlabel metal1 0 1482 34 1516 0 A1
rlabel metal1 0 872 34 906 0 A0
<< end >>
