magic
tech sky130A
magscale 1 2
timestamp 1702568184
<< nwell >>
rect 306 -338 339 -130
rect 0 -425 339 -338
rect 643 -425 721 -130
<< psubdiff >>
rect 237 580 319 604
rect 237 546 262 580
rect 296 546 319 580
rect 237 522 319 546
<< psubdiffcont >>
rect 262 546 296 580
<< poly >>
rect 94 556 193 572
rect 94 522 143 556
rect 177 522 193 556
rect 94 506 193 522
rect 94 479 125 506
rect 262 247 328 258
rect 262 233 278 247
rect 182 213 278 233
rect 312 213 328 247
rect 182 203 328 213
rect 39 160 124 176
rect 39 126 55 160
rect 89 126 124 160
rect 39 110 124 126
rect 94 49 124 110
rect 182 49 212 203
rect 286 133 352 149
rect 432 133 462 179
rect 286 99 302 133
rect 336 99 462 133
rect 286 83 352 99
rect 432 63 462 99
rect 520 174 550 179
rect 520 158 600 174
rect 520 124 550 158
rect 584 124 600 158
rect 520 109 600 124
rect 520 63 550 109
rect 94 -338 212 -302
rect 120 -372 136 -338
rect 170 -372 186 -338
rect 120 -388 186 -372
<< polycont >>
rect 143 522 177 556
rect 278 213 312 247
rect 55 126 89 160
rect 302 99 336 133
rect 550 124 584 158
rect 136 -372 170 -338
<< locali >>
rect 143 556 177 739
rect 237 580 319 604
rect 237 546 262 580
rect 296 546 319 580
rect 237 522 319 546
rect 143 506 177 522
rect 262 213 278 247
rect 312 213 328 247
rect 39 126 55 160
rect 89 126 105 160
rect 386 158 420 201
rect 224 99 302 133
rect 336 99 352 133
rect 386 124 550 158
rect 584 124 600 158
rect 224 27 258 99
rect 386 41 420 124
rect 48 -188 82 -65
rect 224 -188 258 -65
rect 48 -338 82 -280
rect 48 -372 136 -338
rect 170 -372 186 -338
<< viali >>
rect 143 739 177 773
rect 262 546 296 580
rect 278 213 312 247
rect 55 126 89 160
<< metal1 >>
rect 478 929 488 981
rect 540 963 550 981
rect 540 929 835 963
rect 154 841 164 893
rect 216 875 226 893
rect 216 841 835 875
rect 131 773 189 779
rect 12 739 143 773
rect 177 739 856 773
rect 131 733 189 739
rect 729 678 739 690
rect 12 644 739 678
rect 48 453 82 644
rect 237 580 309 644
rect 474 605 508 644
rect 729 638 739 644
rect 791 638 801 690
rect 237 546 262 580
rect 296 546 309 580
rect 237 522 309 546
rect 36 117 46 169
rect 98 117 108 169
rect 136 23 170 285
rect 259 204 269 256
rect 321 204 331 256
rect 562 37 596 205
rect 135 -459 170 -276
rect 318 -363 328 -310
rect 380 -363 390 -310
rect 602 -362 628 -310
rect 680 -362 690 -310
rect 602 -363 690 -362
rect 474 -459 509 -363
rect 729 -949 739 -931
rect 720 -983 739 -949
rect 791 -983 801 -931
<< via1 >>
rect 488 929 540 981
rect 164 841 216 893
rect 739 638 791 690
rect 46 160 98 169
rect 46 126 55 160
rect 55 126 89 160
rect 89 126 98 160
rect 46 117 98 126
rect 269 247 321 256
rect 269 213 278 247
rect 278 213 312 247
rect 312 213 321 247
rect 269 204 321 213
rect 328 -363 380 -310
rect 628 -362 680 -310
rect 739 -983 791 -931
<< metal2 >>
rect 12 719 64 906
rect 164 893 216 1025
rect 488 981 540 1025
rect 488 919 540 929
rect 164 831 216 841
rect 12 685 98 719
rect 46 169 98 685
rect 269 256 321 266
rect 640 256 692 1025
rect 321 204 692 256
rect 739 690 791 700
rect 269 194 321 204
rect 46 107 98 117
rect 328 -310 380 -300
rect 328 -372 380 -363
rect 38 -425 380 -372
rect 628 -310 680 -300
rect 628 -425 680 -362
rect 739 -931 791 638
rect 739 -993 791 -983
use bit_cell  bit_cell_0 ~/Desktop/FabRAM/FE/sram130/bit_cell
timestamp 1702297211
transform 1 0 0 0 1 -1121
box 0 0 720 696
use sky130_fd_pr__nfet_01v8_A6LSUL  m1
timestamp 1702552054
transform -1 0 109 0 1 -19
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_A6LSUL  m2
timestamp 1702552054
transform 1 0 197 0 1 -19
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP#0  m3
timestamp 1702552054
transform -1 0 109 0 1 -234
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP#0  m4
timestamp 1702552054
transform 1 0 197 0 1 -234
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_5YUHNA  m5
timestamp 1702553317
transform -1 0 447 0 1 -163
box -109 -262 109 262
use sky130_fd_pr__nfet_01v8_JB3UY8  m6
timestamp 1702553317
transform -1 0 447 0 1 405
box -73 -226 73 226
use sky130_fd_pr__pfet_01v8_5YUHNA  m7
timestamp 1702553317
transform 1 0 535 0 1 -163
box -109 -262 109 262
use sky130_fd_pr__nfet_01v8_JB3UY8  m8
timestamp 1702553317
transform 1 0 535 0 1 405
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_VJ5ZNR  m9
timestamp 1702559342
transform 1 0 109 0 1 369
box -73 -110 73 110
<< end >>
