magic
tech sky130A
magscale 1 2
timestamp 1702553317
<< error_p >>
rect -239 123 -181 129
rect -239 89 -227 123
rect 97 104 157 142
rect 181 123 239 129
rect 181 89 193 123
rect -239 83 -181 89
rect 181 83 239 89
rect -449 -89 -391 -83
rect -29 -89 29 -83
rect 391 -89 449 -83
rect -449 -123 -437 -89
rect -449 -129 -391 -123
rect -113 -142 -53 -104
rect -29 -123 -17 -89
rect -29 -129 29 -123
rect 307 -142 367 -104
rect 391 -123 403 -89
rect 391 -129 449 -123
<< nwell >>
rect -323 104 -97 142
rect 97 104 323 142
rect -533 -104 533 104
rect -533 -142 -307 -104
rect -113 -142 113 -104
rect 307 -142 533 -104
<< pmos >>
rect -435 -42 -405 42
rect -225 -42 -195 42
rect -15 -42 15 42
rect 195 -42 225 42
rect 405 -42 435 42
<< pdiff >>
rect -497 30 -435 42
rect -497 -30 -485 30
rect -451 -30 -435 30
rect -497 -42 -435 -30
rect -405 30 -343 42
rect -405 -30 -389 30
rect -355 -30 -343 30
rect -405 -42 -343 -30
rect -287 30 -225 42
rect -287 -30 -275 30
rect -241 -30 -225 30
rect -287 -42 -225 -30
rect -195 30 -133 42
rect -195 -30 -179 30
rect -145 -30 -133 30
rect -195 -42 -133 -30
rect -77 30 -15 42
rect -77 -30 -65 30
rect -31 -30 -15 30
rect -77 -42 -15 -30
rect 15 30 77 42
rect 15 -30 31 30
rect 65 -30 77 30
rect 15 -42 77 -30
rect 133 30 195 42
rect 133 -30 145 30
rect 179 -30 195 30
rect 133 -42 195 -30
rect 225 30 287 42
rect 225 -30 241 30
rect 275 -30 287 30
rect 225 -42 287 -30
rect 343 30 405 42
rect 343 -30 355 30
rect 389 -30 405 30
rect 343 -42 405 -30
rect 435 30 497 42
rect 435 -30 451 30
rect 485 -30 497 30
rect 435 -42 497 -30
<< pdiffc >>
rect -485 -30 -451 30
rect -389 -30 -355 30
rect -275 -30 -241 30
rect -179 -30 -145 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 145 -30 179 30
rect 241 -30 275 30
rect 355 -30 389 30
rect 451 -30 485 30
<< poly >>
rect -243 123 -177 139
rect -243 89 -227 123
rect -193 89 -177 123
rect -243 73 -177 89
rect 177 123 243 139
rect 177 89 193 123
rect 227 89 243 123
rect 177 73 243 89
rect -435 42 -405 68
rect -225 42 -195 73
rect -15 42 15 68
rect 195 42 225 73
rect 405 42 435 68
rect -435 -73 -405 -42
rect -225 -68 -195 -42
rect -15 -73 15 -42
rect 195 -68 225 -42
rect 405 -73 435 -42
rect -453 -89 -387 -73
rect -453 -123 -437 -89
rect -403 -123 -387 -89
rect -453 -139 -387 -123
rect -33 -89 33 -73
rect -33 -123 -17 -89
rect 17 -123 33 -89
rect -33 -139 33 -123
rect 387 -89 453 -73
rect 387 -123 403 -89
rect 437 -123 453 -89
rect 387 -139 453 -123
<< polycont >>
rect -227 89 -193 123
rect 193 89 227 123
rect -437 -123 -403 -89
rect -17 -123 17 -89
rect 403 -123 437 -89
<< locali >>
rect -243 89 -227 123
rect -193 89 -177 123
rect 177 89 193 123
rect 227 89 243 123
rect -485 30 -451 46
rect -485 -46 -451 -30
rect -389 30 -355 46
rect -389 -46 -355 -30
rect -275 30 -241 46
rect -275 -46 -241 -30
rect -179 30 -145 46
rect -179 -46 -145 -30
rect -65 30 -31 46
rect -65 -46 -31 -30
rect 31 30 65 46
rect 31 -46 65 -30
rect 145 30 179 46
rect 145 -46 179 -30
rect 241 30 275 46
rect 241 -46 275 -30
rect 355 30 389 46
rect 355 -46 389 -30
rect 451 30 485 46
rect 451 -46 485 -30
rect -453 -123 -437 -89
rect -403 -123 -387 -89
rect -33 -123 -17 -89
rect 17 -123 33 -89
rect 387 -123 403 -89
rect 437 -123 453 -89
<< viali >>
rect -227 89 -193 123
rect 193 89 227 123
rect -485 -30 -451 30
rect -389 -30 -355 30
rect -275 -30 -241 30
rect -179 -30 -145 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 145 -30 179 30
rect 241 -30 275 30
rect 355 -30 389 30
rect 451 -30 485 30
rect -437 -123 -403 -89
rect -17 -123 17 -89
rect 403 -123 437 -89
<< metal1 >>
rect -239 123 -181 129
rect -239 89 -227 123
rect -193 89 -181 123
rect -239 83 -181 89
rect 181 123 239 129
rect 181 89 193 123
rect 227 89 239 123
rect 181 83 239 89
rect -491 30 -445 42
rect -491 -30 -485 30
rect -451 -30 -445 30
rect -491 -42 -445 -30
rect -395 30 -349 42
rect -395 -30 -389 30
rect -355 -30 -349 30
rect -395 -42 -349 -30
rect -281 30 -235 42
rect -281 -30 -275 30
rect -241 -30 -235 30
rect -281 -42 -235 -30
rect -185 30 -139 42
rect -185 -30 -179 30
rect -145 -30 -139 30
rect -185 -42 -139 -30
rect -71 30 -25 42
rect -71 -30 -65 30
rect -31 -30 -25 30
rect -71 -42 -25 -30
rect 25 30 71 42
rect 25 -30 31 30
rect 65 -30 71 30
rect 25 -42 71 -30
rect 139 30 185 42
rect 139 -30 145 30
rect 179 -30 185 30
rect 139 -42 185 -30
rect 235 30 281 42
rect 235 -30 241 30
rect 275 -30 281 30
rect 235 -42 281 -30
rect 349 30 395 42
rect 349 -30 355 30
rect 389 -30 395 30
rect 349 -42 395 -30
rect 445 30 491 42
rect 445 -30 451 30
rect 485 -30 491 30
rect 445 -42 491 -30
rect -449 -89 -391 -83
rect -449 -123 -437 -89
rect -403 -123 -391 -89
rect -449 -129 -391 -123
rect -29 -89 29 -83
rect -29 -123 -17 -89
rect 17 -123 29 -89
rect -29 -129 29 -123
rect 391 -89 449 -83
rect 391 -123 403 -89
rect 437 -123 449 -89
rect 391 -129 449 -123
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 1 nf 5 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
