magic
tech sky130A
magscale 1 2
timestamp 1702392485
<< nwell >>
rect 0 488 330 696
<< nmos >>
rect 206 201 236 285
<< pmos >>
rect 206 550 236 634
<< ndiff >>
rect 148 273 206 285
rect 148 213 160 273
rect 194 213 206 273
rect 148 201 206 213
rect 236 273 294 285
rect 236 213 248 273
rect 282 213 294 273
rect 236 201 294 213
<< pdiff >>
rect 148 622 206 634
rect 148 562 160 622
rect 194 562 206 622
rect 148 550 206 562
rect 236 622 294 634
rect 236 562 248 622
rect 282 562 294 622
rect 236 550 294 562
<< ndiffc >>
rect 160 213 194 273
rect 248 213 282 273
<< pdiffc >>
rect 160 562 194 622
rect 248 562 282 622
<< psubdiff >>
rect 36 273 94 297
rect 36 213 48 273
rect 82 213 94 273
rect 36 189 94 213
<< nsubdiff >>
rect 36 622 94 646
rect 36 562 48 622
rect 82 562 94 622
rect 36 538 94 562
<< psubdiffcont >>
rect 48 213 82 273
<< nsubdiffcont >>
rect 48 562 82 622
<< poly >>
rect 206 634 236 660
rect 206 460 236 550
rect 145 444 236 460
rect 145 410 161 444
rect 195 410 236 444
rect 145 394 236 410
rect 206 285 236 394
rect 206 175 236 201
<< polycont >>
rect 161 410 195 444
<< locali >>
rect 36 622 194 638
rect 36 562 48 622
rect 82 562 160 622
rect 36 546 194 562
rect 248 622 282 638
rect 248 444 282 562
rect 145 410 161 444
rect 195 410 211 444
rect 48 273 194 289
rect 82 213 160 273
rect 48 197 194 213
rect 248 273 282 410
rect 248 197 282 213
<< viali >>
rect 160 562 194 622
rect 248 562 282 622
rect 161 410 195 444
rect 248 410 282 444
rect 160 213 194 273
rect 248 213 282 273
<< metal1 >>
rect 0 662 330 696
rect 160 634 194 662
rect 154 622 200 634
rect 154 562 160 622
rect 194 562 200 622
rect 154 550 200 562
rect 242 622 288 634
rect 242 562 248 622
rect 282 562 288 622
rect 242 550 288 562
rect 149 444 207 450
rect 0 410 161 444
rect 195 410 207 444
rect 149 404 207 410
rect 236 444 294 450
rect 236 410 248 444
rect 282 410 330 444
rect 236 404 294 410
rect 154 273 200 285
rect 154 213 160 273
rect 194 213 200 273
rect 154 201 200 213
rect 242 273 288 285
rect 242 213 248 273
rect 282 213 288 273
rect 242 201 288 213
rect 160 172 194 201
rect 0 138 330 172
<< labels >>
rlabel metal1 296 410 330 444 0 B
rlabel metal1 0 662 34 696 0 VDD
rlabel metal1 0 410 34 444 0 A
rlabel metal1 0 138 34 172 0 VSS
<< end >>
