magic
tech sky130A
magscale 1 2
timestamp 1702826916
<< nwell >>
rect 0 488 394 696
<< pwell >>
rect 10 175 384 311
<< nmos >>
rect 94 201 124 285
rect 182 201 212 285
rect 270 201 300 285
<< pmos >>
rect 94 550 124 634
rect 182 550 212 634
rect 270 550 300 634
<< ndiff >>
rect 36 260 94 285
rect 36 226 48 260
rect 82 226 94 260
rect 36 201 94 226
rect 124 260 182 285
rect 124 226 136 260
rect 170 226 182 260
rect 124 201 182 226
rect 212 260 270 285
rect 212 226 224 260
rect 258 226 270 260
rect 212 201 270 226
rect 300 260 358 285
rect 300 226 312 260
rect 346 226 358 260
rect 300 201 358 226
<< pdiff >>
rect 36 609 94 634
rect 36 575 48 609
rect 82 575 94 609
rect 36 550 94 575
rect 124 609 182 634
rect 124 575 136 609
rect 170 575 182 609
rect 124 550 182 575
rect 212 609 270 634
rect 212 575 224 609
rect 258 575 270 609
rect 212 550 270 575
rect 300 609 358 634
rect 300 575 312 609
rect 346 575 358 609
rect 300 550 358 575
<< ndiffc >>
rect 48 226 82 260
rect 136 226 170 260
rect 224 226 258 260
rect 312 226 346 260
<< pdiffc >>
rect 48 575 82 609
rect 136 575 170 609
rect 224 575 258 609
rect 312 575 346 609
<< poly >>
rect 94 634 124 660
rect 182 634 212 660
rect 270 634 300 660
rect 94 519 124 550
rect 44 503 124 519
rect 44 469 60 503
rect 94 469 124 503
rect 44 453 124 469
rect 94 285 124 453
rect 182 448 212 550
rect 170 432 224 448
rect 170 398 180 432
rect 214 398 224 432
rect 170 382 224 398
rect 182 285 212 382
rect 270 373 300 550
rect 270 357 350 373
rect 270 323 300 357
rect 334 323 350 357
rect 270 307 350 323
rect 270 285 300 307
rect 94 175 124 201
rect 182 175 212 201
rect 270 175 300 201
<< polycont >>
rect 60 469 94 503
rect 180 398 214 432
rect 300 323 334 357
<< locali >>
rect 48 609 82 638
rect 48 546 82 575
rect 136 609 170 638
rect 136 546 170 575
rect 224 609 258 638
rect 224 546 258 575
rect 312 609 346 638
rect 312 546 346 575
rect 44 469 60 503
rect 94 469 110 503
rect 164 398 180 432
rect 214 398 230 432
rect 164 323 180 357
rect 214 323 300 357
rect 334 323 350 357
rect 48 260 82 289
rect 48 197 82 226
rect 136 260 170 289
rect 136 197 170 226
rect 224 260 258 289
rect 224 197 258 226
rect 312 260 346 289
rect 312 197 346 226
<< viali >>
rect 48 575 82 609
rect 136 575 170 609
rect 224 575 258 609
rect 312 575 346 609
rect 60 469 94 503
rect 180 398 214 432
rect 180 323 214 357
rect 48 226 82 260
rect 136 226 170 260
rect 224 226 258 260
rect 312 226 346 260
<< metal1 >>
rect 0 662 394 696
rect 48 634 82 662
rect 224 634 258 662
rect 42 609 88 634
rect 42 575 48 609
rect 82 575 88 609
rect 42 550 88 575
rect 130 609 176 634
rect 130 575 136 609
rect 170 575 176 609
rect 130 550 176 575
rect 218 609 264 634
rect 218 575 224 609
rect 258 575 264 609
rect 218 550 264 575
rect 306 609 352 634
rect 306 575 312 609
rect 346 575 352 609
rect 306 550 352 575
rect 136 522 170 550
rect 312 522 346 550
rect 0 503 106 522
rect 0 488 60 503
rect 48 469 60 488
rect 94 469 106 503
rect 136 488 346 522
rect 48 463 106 469
rect 312 444 346 488
rect 168 432 226 438
rect 0 398 180 432
rect 214 398 226 432
rect 168 392 226 398
rect 312 410 394 444
rect 168 357 226 363
rect 168 351 180 357
rect 0 323 180 351
rect 214 323 226 357
rect 0 317 226 323
rect 312 285 346 410
rect 42 260 88 285
rect 42 226 48 260
rect 82 226 88 260
rect 42 201 88 226
rect 130 260 176 285
rect 130 226 136 260
rect 170 226 176 260
rect 130 201 176 226
rect 218 260 264 285
rect 218 226 224 260
rect 258 226 264 260
rect 218 201 264 226
rect 306 260 352 285
rect 306 226 312 260
rect 346 226 352 260
rect 306 201 352 226
rect 48 172 82 201
rect 0 138 394 172
<< labels >>
flabel metal1 s 0 662 34 696 0 FreeSans 44 0 0 0 VDD
port 1 nsew
flabel metal1 s 0 138 34 172 0 FreeSans 44 0 0 0 VSS
port 2 nsew
flabel metal1 s 360 410 394 444 0 FreeSans 44 0 0 0 Y
port 3 nsew
flabel metal1 s 0 317 34 351 0 FreeSans 44 0 0 0 C
port 4 nsew
flabel metal1 s 0 398 34 432 0 FreeSans 44 0 0 0 B
port 5 nsew
flabel metal1 s 0 488 34 522 0 FreeSans 44 0 0 0 A
port 6 nsew
<< end >>
