magic
tech sky130A
magscale 1 2
timestamp 1702826916
<< nwell >>
rect -166 349 -73 557
<< nmos >>
rect 633 62 663 146
rect 939 62 969 146
rect 1244 62 1274 146
rect 1550 62 1580 146
<< pmos >>
rect 633 411 663 495
rect 939 411 969 495
rect 1244 411 1274 495
rect 1550 411 1580 495
<< ndiff >>
rect 445 134 503 146
rect 445 74 457 134
rect 491 74 503 134
rect 445 62 503 74
rect 751 134 809 146
rect 751 74 763 134
rect 797 74 809 134
rect 751 62 809 74
rect 1056 134 1114 146
rect 1056 74 1068 134
rect 1102 74 1114 134
rect 1056 62 1114 74
rect 1362 134 1420 146
rect 1362 74 1374 134
rect 1408 74 1420 134
rect 1362 62 1420 74
<< pdiff >>
rect 445 483 503 495
rect 445 423 457 483
rect 491 423 503 483
rect 445 411 503 423
rect 751 483 809 495
rect 751 423 763 483
rect 797 423 809 483
rect 751 411 809 423
rect 1056 483 1114 495
rect 1056 423 1068 483
rect 1102 423 1114 483
rect 1056 411 1114 423
rect 1362 483 1420 495
rect 1362 423 1374 483
rect 1408 423 1420 483
rect 1362 411 1420 423
<< ndiffc >>
rect 457 74 491 134
rect 763 74 797 134
rect 1068 74 1102 134
rect 1374 74 1408 134
<< pdiffc >>
rect 457 423 491 483
rect 763 423 797 483
rect 1068 423 1102 483
rect 1374 423 1408 483
<< poly >>
rect 633 495 663 521
rect 939 495 969 521
rect 1244 495 1274 521
rect 1550 495 1580 521
rect -110 305 -44 321
rect 21 305 51 385
rect -110 271 -94 305
rect -60 271 51 305
rect 109 299 139 386
rect -110 255 -44 271
rect 21 172 51 271
rect 93 283 159 299
rect 93 249 109 283
rect 143 249 159 283
rect 93 233 159 249
rect 201 283 255 299
rect 327 283 357 385
rect 201 249 211 283
rect 245 249 357 283
rect 201 233 255 249
rect 109 172 139 233
rect 327 172 357 249
rect 415 172 445 385
rect 507 283 561 299
rect 633 283 663 411
rect 507 249 517 283
rect 551 249 663 283
rect 507 233 561 249
rect 633 146 663 249
rect 721 172 751 385
rect 813 283 867 299
rect 939 283 969 411
rect 813 249 823 283
rect 857 249 969 283
rect 813 233 867 249
rect 939 146 969 249
rect 1026 169 1056 386
rect 1118 283 1172 299
rect 1244 283 1274 411
rect 1118 249 1128 283
rect 1162 249 1274 283
rect 1118 233 1172 249
rect 1244 146 1274 249
rect 1332 172 1362 385
rect 1424 283 1478 299
rect 1550 283 1580 411
rect 1424 249 1434 283
rect 1468 249 1580 283
rect 1424 233 1478 249
rect 1550 146 1580 249
rect 633 36 663 62
rect 939 36 969 62
rect 1244 36 1274 62
rect 1550 36 1580 62
<< polycont >>
rect -94 271 -60 305
rect 109 249 143 283
rect 211 249 245 283
rect 517 249 551 283
rect 823 249 857 283
rect 1128 249 1162 283
rect 1434 249 1468 283
<< locali >>
rect 457 483 491 499
rect 159 407 245 441
rect 763 483 797 499
rect 491 423 551 441
rect 457 407 551 423
rect 1068 483 1102 499
rect 797 423 857 441
rect 763 407 857 423
rect 1374 483 1408 499
rect 1102 423 1162 441
rect 1068 407 1162 423
rect 1408 423 1468 441
rect 1374 407 1468 423
rect -94 305 -60 321
rect -94 255 -60 271
rect -25 283 9 407
rect 211 283 245 407
rect -25 249 109 283
rect 143 249 159 283
rect -25 150 9 249
rect 211 150 245 249
rect 281 150 315 407
rect 517 283 551 407
rect 517 150 551 249
rect 587 150 621 407
rect 823 283 857 407
rect 823 150 857 249
rect 892 150 926 407
rect 1128 283 1162 407
rect 1128 150 1162 249
rect 1198 150 1232 407
rect 1434 283 1468 407
rect 1434 150 1468 249
rect 1592 218 1626 407
rect 1592 150 1626 184
rect 159 116 245 150
rect 457 134 551 150
rect 491 116 551 134
rect 763 134 857 150
rect 457 58 491 74
rect 797 116 857 134
rect 1068 134 1162 150
rect 763 58 797 74
rect 1102 116 1162 134
rect 1374 134 1468 150
rect 1068 58 1102 74
rect 1408 116 1468 134
rect 1374 58 1408 74
<< viali >>
rect 457 423 491 483
rect 763 423 797 483
rect 1068 423 1102 483
rect 1374 423 1408 483
rect -94 271 -60 305
rect 1592 184 1626 218
rect 457 74 491 134
rect 763 74 797 134
rect 1068 74 1102 134
rect 1374 74 1408 134
<< metal1 >>
rect -166 523 1674 557
rect 63 495 97 523
rect 369 495 403 523
rect 674 495 708 523
rect 980 495 1014 523
rect 1286 495 1320 523
rect 1504 495 1538 523
rect 451 483 497 495
rect 451 423 457 483
rect 491 423 497 483
rect 451 411 497 423
rect 757 483 803 495
rect 757 423 763 483
rect 797 423 803 483
rect 757 411 803 423
rect 1062 483 1108 495
rect 1062 423 1068 483
rect 1102 423 1108 483
rect 1062 411 1108 423
rect 1368 483 1414 495
rect 1368 423 1374 483
rect 1408 423 1414 483
rect 1368 411 1414 423
rect 139 329 1674 363
rect -106 305 -48 311
rect 139 305 167 329
rect -166 271 -94 305
rect -60 271 167 305
rect -106 265 -48 271
rect 1580 218 1638 224
rect 1580 184 1592 218
rect 1626 184 1674 218
rect 1580 178 1638 184
rect 451 134 497 146
rect 451 74 457 134
rect 491 74 497 134
rect 451 62 497 74
rect 757 134 803 146
rect 757 74 763 134
rect 797 74 803 134
rect 757 62 803 74
rect 1062 134 1108 146
rect 1062 74 1068 134
rect 1102 74 1108 134
rect 1062 62 1108 74
rect 1368 134 1414 146
rect 1368 74 1374 134
rect 1408 74 1414 134
rect 1368 62 1414 74
rect 63 33 97 62
rect 369 33 403 62
rect 675 33 709 62
rect 980 33 1014 62
rect 1504 33 1538 62
rect -166 -1 1674 33
use sky130_fd_pr__nfet_01v8_A6LSUL  m1
timestamp 1702809544
transform -1 0 36 0 1 104
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_A6LSUL  m2
timestamp 1702809544
transform 1 0 124 0 1 104
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_A6LSUL  m3
timestamp 1702809544
transform -1 0 342 0 1 104
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_A6LSUL  m4
timestamp 1702809544
transform 1 0 430 0 1 104
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_A6LSUL  m5
timestamp 1702809544
transform -1 0 648 0 1 104
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_A6LSUL  m6
timestamp 1702809544
transform 1 0 736 0 1 104
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_A6LSUL  m7
timestamp 1702809544
transform -1 0 953 0 1 104
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_A6LSUL  m8
timestamp 1702809544
transform 1 0 1041 0 1 104
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_A6LSUL  m9
timestamp 1702809544
transform -1 0 1259 0 1 104
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_A6LSUL  m10
timestamp 1702809544
transform -1 0 1347 0 1 104
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_A6LSUL  m11
timestamp 1702809544
transform 1 0 1565 0 1 104
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m12
timestamp 1702809649
transform -1 0 36 0 1 453
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m13
timestamp 1702809649
transform 1 0 124 0 1 453
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m14
timestamp 1702809649
transform -1 0 342 0 1 453
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m15
timestamp 1702809649
transform 1 0 430 0 1 453
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m16
timestamp 1702809649
transform -1 0 648 0 1 453
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m17
timestamp 1702809649
transform 1 0 736 0 1 453
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m18
timestamp 1702809649
transform -1 0 953 0 1 453
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m19
timestamp 1702809649
transform 1 0 1041 0 1 453
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m20
timestamp 1702809649
transform -1 0 1259 0 1 453
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m21
timestamp 1702809649
transform 1 0 1347 0 1 453
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m22
timestamp 1702809649
transform 1 0 1565 0 1 453
box -109 -104 109 104
use nand2_f  nand2_f_0 ~/Desktop/FabRAM/FE/sram130/nand2
timestamp 1702826916
transform 1 0 1674 0 1 -139
box 0 138 306 696
use not_f  not_f_0 ~/Desktop/FabRAM/FE/sram130/not
timestamp 1702826916
transform 1 0 1980 0 1 -139
box 0 138 330 696
<< end >>
