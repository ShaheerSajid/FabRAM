.title characterizer
.include /home/shaheer/Desktop/FabRAM/FE/out/sram1024x32.spi
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

      .tran 0.01179285n 23.585700000000003n 11.792850000000001n
      .control
      set hcopydevtype = svg
      run
      meas tran tdiff_cell_rise TRIG v(clk) VAL=0.9 RISE=1 TARG v(Q0) VAL=0.9 RISE=1 
      meas tran tdiff_tran_rise TRIG v(Q0)  VAL=0.18000000000000002 RISE=1 TARG v(Q0) VAL=1.62 RISE=1 
      meas tran tdiff_cell_fall TRIG v(clk) VAL=0.9 RISE=2 TARG v(Q0) VAL=0.9 FALL=1 
      meas tran tdiff_tran_fall TRIG v(Q0)  VAL=1.62 FALL=1 TARG v(Q0) VAL=0.18000000000000002 FALL=1 

      echo "$&tdiff_cell_rise,$&tdiff_tran_rise $&tdiff_cell_fall,$&tdiff_tran_fall" > log/sim_0.35857_0.03432.text
      hardcopy log/sim_0.35857_0.03432.svg v(clk)+9.0 v(Q0)+7.2 v(x0.PCHG)+5.4 v(x0.WLEN)+3.6 v(x0.SAEN)+1.8 v(x0.WREN) v(x0.x8.RBL)
      exit
      .endc
      
Vpower VDD 0 1.8
Vgnd VSS 0 0
Vclk clk VSS DC 0V PULSE(0V 1.8V 0ns 0.44821249999999996ns 0.44821249999999996ns 2.5ns 5.896425000000001ns)
Vaddr addr VSS DC 0V PULSE(0V 1.8V 0s 1ps 1ps 2.5ns 11.792850000000001ns)
Vdin din VSS DC 0V PULSE(0V 1.8V 0s 1ps 1ps 2.5ns 11.792850000000001ns)
Vwrite write VSS DC 0V PULSE(0V 1.8V 0s 1ps 1ps 11.792850000000001ns 23.585700000000003ns)
X0 VDD VSS clk addr addr addr addr addr addr addr addr addr addr din din din din din din din din din din din din din din din din din din din din din din din din din din din din din din din din Q0 Q1 Q2 Q3 Q4 Q5 Q6 Q7 Q8 Q9 Q10 Q11 Q12 Q13 Q14 Q15 Q16 Q17 Q18 Q19 Q20 Q21 Q22 Q23 Q24 Q25 Q26 Q27 Q28 Q29 Q30 Q31 write VDD sram1024x32
C0 Q0 VSS 0.03432p
