magic
tech sky130A
magscale 1 2
timestamp 1702809649
<< nwell >>
rect 658 -841 798 -633
<< ndiff >>
rect 3148 -476 3206 -464
rect 3148 -612 3160 -476
rect 3194 -612 3206 -476
rect 3148 -624 3206 -612
<< pdiff >>
rect 3148 -102 3206 -90
rect 3148 -238 3160 -102
rect 3194 -238 3206 -102
rect 3148 -250 3206 -238
<< ndiffc >>
rect 3160 -612 3194 -476
<< pdiffc >>
rect 3160 -238 3194 -102
<< poly >>
rect 2884 -9 2950 7
rect 2884 -43 2900 -9
rect 2934 -43 2950 -9
rect 2884 -59 2950 -43
rect 2900 -64 2930 -59
rect 3118 -342 3148 -276
rect 3336 -342 3366 -250
rect 2850 -358 2930 -342
rect 2850 -392 2866 -358
rect 2900 -392 2930 -358
rect 2850 -408 2930 -392
rect 3057 -358 3148 -342
rect 3057 -392 3073 -358
rect 3107 -392 3148 -358
rect 3057 -408 3148 -392
rect 3275 -358 3366 -342
rect 3275 -392 3291 -358
rect 3325 -392 3366 -358
rect 3520 -324 3586 -308
rect 3520 -358 3536 -324
rect 3570 -358 3586 -324
rect 3520 -374 3586 -358
rect 3275 -408 3366 -392
rect 2900 -438 2930 -408
rect 3118 -438 3148 -408
rect 3336 -464 3366 -408
rect 3547 -438 3577 -374
<< polycont >>
rect 2900 -43 2934 -9
rect 2866 -392 2900 -358
rect 3073 -392 3107 -358
rect 3291 -392 3325 -358
rect 3536 -358 3570 -324
<< locali >>
rect 3054 -9 3088 60
rect 2884 -43 2900 -9
rect 2934 -43 3570 -9
rect 3160 -102 3194 -86
rect 2866 -358 2900 -342
rect 2866 -408 2900 -392
rect 2942 -358 2976 -254
rect 3160 -358 3194 -238
rect 2942 -392 3073 -358
rect 3107 -392 3123 -358
rect 3160 -392 3291 -358
rect 3325 -392 3341 -358
rect 2942 -460 2976 -392
rect 3160 -476 3194 -392
rect 3378 -430 3412 -254
rect 3536 -324 3570 -43
rect 3536 -374 3570 -358
rect 3378 -460 3535 -430
rect 3412 -464 3535 -460
rect 3160 -716 3194 -612
rect 3049 -750 3194 -716
rect 3049 -954 3083 -750
rect 3049 -988 3128 -954
<< viali >>
rect 3160 -238 3194 -102
rect 2866 -392 2900 -358
rect 3160 -612 3194 -476
<< metal1 >>
rect -93 272 34 306
rect -93 -280 -59 272
rect 2854 -28 3024 -27
rect 2806 -62 3461 -28
rect 2854 -90 2888 -62
rect 3072 -90 3106 -62
rect 3154 -102 3200 -90
rect 3154 -238 3160 -102
rect 3194 -238 3200 -102
rect 3290 -166 3324 -62
rect 3154 -250 3200 -238
rect -155 -314 391 -280
rect 2806 -314 2900 -280
rect 2866 -352 2900 -314
rect 2854 -358 2912 -352
rect 2854 -392 2866 -358
rect 2900 -392 3623 -358
rect 2854 -398 2912 -392
rect 3589 -464 3623 -392
rect 3154 -476 3200 -464
rect 2806 -586 2848 -552
rect 2849 -586 2854 -552
rect 3154 -612 3160 -476
rect 3194 -612 3200 -476
rect 3154 -624 3200 -612
rect 658 -667 798 -633
rect 2854 -653 2888 -624
rect 3072 -653 3106 -624
rect 3290 -653 3324 -548
rect 772 -861 806 -667
rect 2854 -687 3449 -653
rect 622 -885 624 -879
rect 658 -919 738 -885
rect 704 -972 738 -919
rect 704 -1006 798 -972
rect 658 -1191 798 -1157
use del_cell  del_cell_0
timestamp 1702809649
transform 1 0 496 0 1 1
box -166 -1 2310 557
use del_cell  del_cell_1
timestamp 1702809649
transform 1 0 496 0 1 -585
box -166 -1 2310 557
use sky130_fd_pr__nfet_01v8_BBXUYH  m1
timestamp 1702809544
transform 1 0 2915 0 1 -544
box -73 -106 73 106
use sky130_fd_pr__pfet_01v8_5C6TXA  m2
timestamp 1702809544
transform 1 0 2915 0 1 -170
box -109 -142 109 142
use sky130_fd_pr__pfet_01v8_5C6TXA  m3
timestamp 1702809544
transform 1 0 3133 0 1 -170
box -109 -142 109 142
use sky130_fd_pr__nfet_01v8_BBXUYH  m4
timestamp 1702809544
transform 1 0 3133 0 1 -544
box -73 -106 73 106
use sky130_fd_pr__pfet_01v8_4Y88KP  m5
timestamp 1702809649
transform 1 0 3351 0 1 -208
box -109 -104 109 104
use sky130_fd_pr__nfet_01v8_A6LSUL  m6
timestamp 1702809544
transform 1 0 3351 0 1 -506
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_BBXUYH  m7
timestamp 1702809544
transform 1 0 3562 0 1 -544
box -73 -106 73 106
use sky130_fd_pr__pfet_01v8_4Y88KP  m8
timestamp 1702809649
transform 1 0 1485 0 1 -738
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m9
timestamp 1702809649
transform 1 0 1703 0 1 -738
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m10
timestamp 1702809649
transform 1 0 1595 0 1 -946
box -109 -104 109 104
use nand2_f  nand2_f_0 ~/Desktop/FabRAM/FE/sram130/nand2
timestamp 1702393006
transform 1 0 3083 0 1 -1456
box 0 138 306 696
use nand2_f  nand2_f_1
timestamp 1702393006
transform 1 0 798 0 1 -1329
box 0 138 306 696
use not_f  not_f_0 ~/Desktop/FabRAM/FE/sram130/not
timestamp 1702392485
transform 1 0 0 0 1 -138
box 0 138 330 696
use not_f  not_f_1
timestamp 1702392485
transform 1 0 2806 0 1 -137
box 0 138 330 696
use not_f  not_f_2
timestamp 1702392485
transform 1 0 3389 0 1 -1456
box 0 138 330 696
use not_f  not_f_3
timestamp 1702392485
transform 1 0 328 0 1 -1329
box 0 138 330 696
<< end >>
