magic
tech sky130A
magscale 1 2
timestamp 1703823919
<< nwell >>
rect 428 1184 1304 1392
rect 99 488 1304 696
<< pwell >>
rect 438 871 1294 1007
rect 109 311 219 323
rect 109 175 419 311
rect 438 175 1294 311
rect 109 163 219 175
<< nmos >>
rect 522 897 552 981
rect 610 897 640 981
rect 828 897 858 981
rect 916 897 946 981
rect 1004 897 1034 981
rect 1092 897 1122 981
rect 1180 897 1210 981
rect 305 201 335 285
rect 522 201 552 285
rect 610 201 640 285
rect 828 201 858 285
rect 916 201 946 285
rect 1004 201 1034 285
rect 1092 201 1122 285
rect 1180 201 1210 285
<< pmos >>
rect 522 1246 552 1330
rect 610 1246 640 1330
rect 828 1246 858 1330
rect 916 1246 946 1330
rect 1004 1246 1034 1330
rect 1092 1246 1122 1330
rect 1180 1246 1210 1330
rect 305 550 335 634
rect 522 550 552 634
rect 610 550 640 634
rect 828 550 858 634
rect 916 550 946 634
rect 1004 550 1034 634
rect 1092 550 1122 634
rect 1180 550 1210 634
<< ndiff >>
rect 464 956 522 981
rect 464 922 476 956
rect 510 922 522 956
rect 464 897 522 922
rect 552 956 610 981
rect 552 922 564 956
rect 598 922 610 956
rect 552 897 610 922
rect 640 956 698 981
rect 640 922 652 956
rect 686 922 698 956
rect 640 897 698 922
rect 770 956 828 981
rect 770 922 782 956
rect 816 922 828 956
rect 770 897 828 922
rect 858 956 916 981
rect 858 922 870 956
rect 904 922 916 956
rect 858 897 916 922
rect 946 956 1004 981
rect 946 922 958 956
rect 992 922 1004 956
rect 946 897 1004 922
rect 1034 956 1092 981
rect 1034 922 1046 956
rect 1080 922 1092 956
rect 1034 897 1092 922
rect 1122 956 1180 981
rect 1122 922 1134 956
rect 1168 922 1180 956
rect 1122 897 1180 922
rect 1210 956 1268 981
rect 1210 922 1222 956
rect 1256 922 1268 956
rect 1210 897 1268 922
rect 247 260 305 285
rect 247 226 259 260
rect 293 226 305 260
rect 247 201 305 226
rect 335 260 393 285
rect 335 226 347 260
rect 381 226 393 260
rect 335 201 393 226
rect 464 260 522 285
rect 464 226 476 260
rect 510 226 522 260
rect 464 201 522 226
rect 552 260 610 285
rect 552 226 564 260
rect 598 226 610 260
rect 552 201 610 226
rect 640 260 698 285
rect 640 226 652 260
rect 686 226 698 260
rect 640 201 698 226
rect 770 260 828 285
rect 770 226 782 260
rect 816 226 828 260
rect 770 201 828 226
rect 858 260 916 285
rect 858 226 870 260
rect 904 226 916 260
rect 858 201 916 226
rect 946 260 1004 285
rect 946 226 958 260
rect 992 226 1004 260
rect 946 201 1004 226
rect 1034 260 1092 285
rect 1034 226 1046 260
rect 1080 226 1092 260
rect 1034 201 1092 226
rect 1122 260 1180 285
rect 1122 226 1134 260
rect 1168 226 1180 260
rect 1122 201 1180 226
rect 1210 260 1268 285
rect 1210 226 1222 260
rect 1256 226 1268 260
rect 1210 201 1268 226
<< pdiff >>
rect 464 1305 522 1330
rect 464 1271 476 1305
rect 510 1271 522 1305
rect 464 1246 522 1271
rect 552 1305 610 1330
rect 552 1271 564 1305
rect 598 1271 610 1305
rect 552 1246 610 1271
rect 640 1305 698 1330
rect 640 1271 652 1305
rect 686 1271 698 1305
rect 640 1246 698 1271
rect 770 1305 828 1330
rect 770 1271 782 1305
rect 816 1271 828 1305
rect 770 1246 828 1271
rect 858 1305 916 1330
rect 858 1271 870 1305
rect 904 1271 916 1305
rect 858 1246 916 1271
rect 946 1305 1004 1330
rect 946 1271 958 1305
rect 992 1271 1004 1305
rect 946 1246 1004 1271
rect 1034 1305 1092 1330
rect 1034 1271 1046 1305
rect 1080 1271 1092 1305
rect 1034 1246 1092 1271
rect 1122 1305 1180 1330
rect 1122 1271 1134 1305
rect 1168 1271 1180 1305
rect 1122 1246 1180 1271
rect 1210 1305 1268 1330
rect 1210 1271 1222 1305
rect 1256 1271 1268 1305
rect 1210 1246 1268 1271
rect 247 609 305 634
rect 247 575 259 609
rect 293 575 305 609
rect 247 550 305 575
rect 335 609 393 634
rect 335 575 347 609
rect 381 575 393 609
rect 335 550 393 575
rect 464 609 522 634
rect 464 575 476 609
rect 510 575 522 609
rect 464 550 522 575
rect 552 609 610 634
rect 552 575 564 609
rect 598 575 610 609
rect 552 550 610 575
rect 640 609 698 634
rect 640 575 652 609
rect 686 575 698 609
rect 640 550 698 575
rect 770 609 828 634
rect 770 575 782 609
rect 816 575 828 609
rect 770 550 828 575
rect 858 609 916 634
rect 858 575 870 609
rect 904 575 916 609
rect 858 550 916 575
rect 946 609 1004 634
rect 946 575 958 609
rect 992 575 1004 609
rect 946 550 1004 575
rect 1034 609 1092 634
rect 1034 575 1046 609
rect 1080 575 1092 609
rect 1034 550 1092 575
rect 1122 609 1180 634
rect 1122 575 1134 609
rect 1168 575 1180 609
rect 1122 550 1180 575
rect 1210 609 1268 634
rect 1210 575 1222 609
rect 1256 575 1268 609
rect 1210 550 1268 575
<< ndiffc >>
rect 476 922 510 956
rect 564 922 598 956
rect 652 922 686 956
rect 782 922 816 956
rect 870 922 904 956
rect 958 922 992 956
rect 1046 922 1080 956
rect 1134 922 1168 956
rect 1222 922 1256 956
rect 259 226 293 260
rect 347 226 381 260
rect 476 226 510 260
rect 564 226 598 260
rect 652 226 686 260
rect 782 226 816 260
rect 870 226 904 260
rect 958 226 992 260
rect 1046 226 1080 260
rect 1134 226 1168 260
rect 1222 226 1256 260
<< pdiffc >>
rect 476 1271 510 1305
rect 564 1271 598 1305
rect 652 1271 686 1305
rect 782 1271 816 1305
rect 870 1271 904 1305
rect 958 1271 992 1305
rect 1046 1271 1080 1305
rect 1134 1271 1168 1305
rect 1222 1271 1256 1305
rect 259 575 293 609
rect 347 575 381 609
rect 476 575 510 609
rect 564 575 598 609
rect 652 575 686 609
rect 782 575 816 609
rect 870 575 904 609
rect 958 575 992 609
rect 1046 575 1080 609
rect 1134 575 1168 609
rect 1222 575 1256 609
<< psubdiff >>
rect 135 260 193 297
rect 135 226 147 260
rect 181 226 193 260
rect 135 189 193 226
<< nsubdiff >>
rect 135 609 193 646
rect 135 575 147 609
rect 181 575 193 609
rect 135 538 193 575
<< psubdiffcont >>
rect 147 226 181 260
<< nsubdiffcont >>
rect 147 575 181 609
<< poly >>
rect 522 1330 552 1356
rect 610 1330 640 1356
rect 828 1330 858 1356
rect 916 1330 946 1356
rect 1004 1330 1034 1356
rect 1092 1330 1122 1356
rect 1180 1330 1210 1356
rect 522 1214 552 1246
rect 472 1198 552 1214
rect 472 1164 488 1198
rect 522 1164 552 1198
rect 472 1148 552 1164
rect 522 981 552 1148
rect 610 1069 640 1246
rect 828 1158 858 1246
rect 775 1140 858 1158
rect 916 1140 946 1246
rect 1004 1140 1034 1246
rect 1092 1140 1122 1246
rect 1180 1140 1210 1246
rect 775 1106 785 1140
rect 819 1106 1210 1140
rect 775 1090 858 1106
rect 610 1053 690 1069
rect 610 1019 640 1053
rect 674 1019 690 1053
rect 610 1003 690 1019
rect 610 981 640 1003
rect 828 981 858 1090
rect 916 981 946 1106
rect 1004 981 1034 1106
rect 1092 981 1122 1106
rect 1180 981 1210 1106
rect 522 871 552 897
rect 610 871 640 897
rect 828 871 858 897
rect 916 871 946 897
rect 1004 871 1034 897
rect 1092 871 1122 897
rect 1180 871 1210 897
rect 305 634 335 660
rect 522 634 552 660
rect 610 634 640 660
rect 828 634 858 660
rect 916 634 946 660
rect 1004 634 1034 660
rect 1092 634 1122 660
rect 1180 634 1210 660
rect 305 460 335 550
rect 522 518 552 550
rect 244 444 335 460
rect 472 502 552 518
rect 472 468 488 502
rect 522 468 552 502
rect 472 452 552 468
rect 244 410 260 444
rect 294 410 335 444
rect 244 394 335 410
rect 305 285 335 394
rect 522 285 552 452
rect 610 373 640 550
rect 828 462 858 550
rect 775 444 858 462
rect 916 444 946 550
rect 1004 444 1034 550
rect 1092 444 1122 550
rect 1180 444 1210 550
rect 775 410 785 444
rect 819 410 1210 444
rect 775 394 858 410
rect 610 357 690 373
rect 610 323 640 357
rect 674 323 690 357
rect 610 307 690 323
rect 610 285 640 307
rect 828 285 858 394
rect 916 285 946 410
rect 1004 285 1034 410
rect 1092 285 1122 410
rect 1180 285 1210 410
rect 305 175 335 201
rect 522 175 552 201
rect 610 175 640 201
rect 828 175 858 201
rect 916 175 946 201
rect 1004 175 1034 201
rect 1092 175 1122 201
rect 1180 175 1210 201
<< polycont >>
rect 488 1164 522 1198
rect 785 1106 819 1140
rect 640 1019 674 1053
rect 488 468 522 502
rect 260 410 294 444
rect 785 410 819 444
rect 640 323 674 357
<< locali >>
rect 476 1305 510 1334
rect 476 1242 510 1271
rect 564 1305 598 1334
rect 564 1242 598 1271
rect 652 1305 686 1334
rect 652 1242 686 1271
rect 782 1305 816 1334
rect 782 1242 816 1271
rect 870 1305 904 1334
rect 472 1164 488 1198
rect 522 1164 538 1198
rect 870 1192 904 1271
rect 958 1305 992 1334
rect 958 1242 992 1271
rect 1046 1305 1080 1334
rect 1046 1192 1080 1271
rect 1134 1305 1168 1334
rect 1134 1242 1168 1271
rect 1222 1305 1256 1334
rect 1222 1192 1256 1271
rect 870 1157 1256 1192
rect 1222 1140 1256 1157
rect 768 1106 785 1140
rect 819 1106 835 1140
rect 1222 1054 1256 1106
rect 476 1019 488 1053
rect 522 1019 640 1053
rect 674 1019 690 1053
rect 870 1019 1256 1054
rect 476 956 510 985
rect 476 893 510 922
rect 564 956 598 985
rect 564 893 598 922
rect 652 956 686 985
rect 652 893 686 922
rect 782 956 816 985
rect 782 893 816 922
rect 870 956 904 1019
rect 870 893 904 922
rect 958 956 992 985
rect 958 893 992 922
rect 1046 956 1080 1019
rect 1046 893 1080 922
rect 1134 956 1168 985
rect 1134 893 1168 922
rect 1222 956 1256 1019
rect 1222 893 1256 922
rect 135 609 293 638
rect 135 575 147 609
rect 181 575 259 609
rect 135 546 293 575
rect 347 609 381 638
rect 347 444 381 575
rect 476 609 510 638
rect 476 546 510 575
rect 564 609 598 638
rect 564 546 598 575
rect 652 609 686 638
rect 652 546 686 575
rect 782 609 816 638
rect 782 546 816 575
rect 870 609 904 638
rect 472 468 488 502
rect 522 468 538 502
rect 870 496 904 575
rect 958 609 992 638
rect 958 546 992 575
rect 1046 609 1080 638
rect 1046 496 1080 575
rect 1134 609 1168 638
rect 1134 546 1168 575
rect 1222 609 1256 638
rect 1222 496 1256 575
rect 870 461 1256 496
rect 1222 444 1256 461
rect 244 410 260 444
rect 294 410 310 444
rect 768 410 785 444
rect 819 410 835 444
rect 147 260 293 289
rect 181 226 259 260
rect 147 197 293 226
rect 347 260 381 410
rect 1222 358 1256 410
rect 476 323 488 357
rect 522 323 640 357
rect 674 323 690 357
rect 870 323 1256 358
rect 347 197 381 226
rect 476 260 510 289
rect 476 197 510 226
rect 564 260 598 289
rect 564 197 598 226
rect 652 260 686 289
rect 652 197 686 226
rect 782 260 816 289
rect 782 197 816 226
rect 870 260 904 323
rect 870 197 904 226
rect 958 260 992 289
rect 958 197 992 226
rect 1046 260 1080 323
rect 1046 197 1080 226
rect 1134 260 1168 289
rect 1134 197 1168 226
rect 1222 260 1256 323
rect 1222 197 1256 226
<< viali >>
rect 476 1271 510 1305
rect 564 1271 598 1305
rect 652 1271 686 1305
rect 782 1271 816 1305
rect 870 1271 904 1305
rect 488 1164 522 1198
rect 958 1271 992 1305
rect 1046 1271 1080 1305
rect 1134 1271 1168 1305
rect 1222 1271 1256 1305
rect 785 1106 819 1140
rect 1222 1106 1256 1140
rect 488 1019 522 1053
rect 476 922 510 956
rect 564 922 598 956
rect 652 922 686 956
rect 782 922 816 956
rect 870 922 904 956
rect 958 922 992 956
rect 1046 922 1080 956
rect 1134 922 1168 956
rect 1222 922 1256 956
rect 259 575 293 609
rect 347 575 381 609
rect 476 575 510 609
rect 564 575 598 609
rect 652 575 686 609
rect 782 575 816 609
rect 870 575 904 609
rect 488 468 522 502
rect 958 575 992 609
rect 1046 575 1080 609
rect 1134 575 1168 609
rect 1222 575 1256 609
rect 260 410 294 444
rect 347 410 381 444
rect 785 410 819 444
rect 1222 410 1256 444
rect 259 226 293 260
rect 488 323 522 357
rect 347 226 381 260
rect 476 226 510 260
rect 564 226 598 260
rect 652 226 686 260
rect 782 226 816 260
rect 870 226 904 260
rect 958 226 992 260
rect 1046 226 1080 260
rect 1134 226 1168 260
rect 1222 226 1256 260
<< metal1 >>
rect 0 1358 1304 1392
rect 476 1330 510 1358
rect 652 1330 686 1358
rect 782 1330 816 1358
rect 958 1330 992 1358
rect 1134 1330 1168 1358
rect 470 1305 516 1330
rect 470 1271 476 1305
rect 510 1271 516 1305
rect 470 1246 516 1271
rect 558 1305 604 1330
rect 558 1271 564 1305
rect 598 1271 604 1305
rect 558 1246 604 1271
rect 646 1305 692 1330
rect 646 1271 652 1305
rect 686 1271 692 1305
rect 646 1246 692 1271
rect 776 1305 822 1330
rect 776 1271 782 1305
rect 816 1271 822 1305
rect 776 1246 822 1271
rect 864 1305 910 1330
rect 864 1271 870 1305
rect 904 1271 910 1305
rect 864 1246 910 1271
rect 952 1305 998 1330
rect 952 1271 958 1305
rect 992 1271 998 1305
rect 952 1246 998 1271
rect 1040 1305 1086 1330
rect 1040 1271 1046 1305
rect 1080 1271 1086 1305
rect 1040 1246 1086 1271
rect 1128 1305 1174 1330
rect 1128 1271 1134 1305
rect 1168 1271 1174 1305
rect 1128 1246 1174 1271
rect 1216 1305 1262 1330
rect 1216 1271 1222 1305
rect 1256 1271 1262 1305
rect 1216 1246 1262 1271
rect 476 1198 534 1204
rect 428 1164 488 1198
rect 522 1164 534 1198
rect 428 1158 534 1164
rect 428 1140 462 1158
rect 0 1106 99 1140
rect 89 1088 99 1106
rect 151 1106 462 1140
rect 564 1140 598 1246
rect 773 1140 831 1146
rect 564 1106 785 1140
rect 819 1106 831 1140
rect 151 1088 161 1106
rect 463 1010 473 1062
rect 525 1010 535 1062
rect 652 981 686 1106
rect 773 1100 831 1106
rect 1210 1140 1268 1146
rect 1458 1140 1468 1162
rect 1210 1106 1222 1140
rect 1256 1106 1468 1140
rect 1524 1106 1534 1162
rect 1210 1100 1268 1106
rect 470 956 516 981
rect 470 922 476 956
rect 510 922 516 956
rect 470 897 516 922
rect 558 956 604 981
rect 558 922 564 956
rect 598 922 604 956
rect 558 897 604 922
rect 646 956 692 981
rect 646 922 652 956
rect 686 922 692 956
rect 646 897 692 922
rect 776 956 822 981
rect 776 922 782 956
rect 816 922 822 956
rect 776 897 822 922
rect 864 956 910 981
rect 864 922 870 956
rect 904 922 910 956
rect 864 897 910 922
rect 952 956 998 981
rect 952 922 958 956
rect 992 922 998 956
rect 952 897 998 922
rect 1040 956 1086 981
rect 1040 922 1046 956
rect 1080 922 1086 956
rect 1040 897 1086 922
rect 1128 956 1174 981
rect 1128 922 1134 956
rect 1168 922 1174 956
rect 1128 897 1174 922
rect 1216 956 1262 981
rect 1216 922 1222 956
rect 1256 922 1262 956
rect 1216 897 1262 922
rect 476 868 510 897
rect 782 868 816 897
rect 958 868 992 897
rect 1134 868 1168 897
rect 0 834 1304 868
rect 99 662 1304 696
rect 259 634 293 662
rect 476 634 510 662
rect 652 634 686 662
rect 782 634 816 662
rect 958 634 992 662
rect 1134 634 1168 662
rect 253 609 299 634
rect 253 575 259 609
rect 293 575 299 609
rect 253 550 299 575
rect 341 609 387 634
rect 341 575 347 609
rect 381 575 387 609
rect 341 550 387 575
rect 470 609 516 634
rect 470 575 476 609
rect 510 575 516 609
rect 470 550 516 575
rect 558 609 604 634
rect 558 575 564 609
rect 598 575 604 609
rect 558 550 604 575
rect 646 609 692 634
rect 646 575 652 609
rect 686 575 692 609
rect 646 550 692 575
rect 776 609 822 634
rect 776 575 782 609
rect 816 575 822 609
rect 776 550 822 575
rect 864 609 910 634
rect 864 575 870 609
rect 904 575 910 609
rect 864 550 910 575
rect 952 609 998 634
rect 952 575 958 609
rect 992 575 998 609
rect 952 550 998 575
rect 1040 609 1086 634
rect 1040 575 1046 609
rect 1080 575 1086 609
rect 1040 550 1086 575
rect 1128 609 1174 634
rect 1128 575 1134 609
rect 1168 575 1174 609
rect 1128 550 1174 575
rect 1216 609 1262 634
rect 1216 575 1222 609
rect 1256 575 1262 609
rect 1216 550 1262 575
rect 476 502 534 508
rect 428 468 488 502
rect 522 468 534 502
rect 428 462 534 468
rect 89 410 99 462
rect 151 444 161 462
rect 248 444 306 450
rect 151 410 260 444
rect 294 410 306 444
rect 248 404 306 410
rect 335 444 393 450
rect 428 444 462 462
rect 335 410 347 444
rect 381 410 462 444
rect 564 444 598 550
rect 773 444 831 450
rect 564 410 785 444
rect 819 410 831 444
rect 335 404 393 410
rect 463 314 473 366
rect 525 314 535 366
rect 652 285 686 410
rect 773 404 831 410
rect 1210 444 1268 450
rect 1552 444 1562 466
rect 1210 410 1222 444
rect 1256 410 1562 444
rect 1618 410 1628 466
rect 1210 404 1268 410
rect 2652 369 2686 1499
rect 2652 334 2774 369
rect 253 260 299 285
rect 253 226 259 260
rect 293 226 299 260
rect 253 201 299 226
rect 341 260 387 285
rect 341 226 347 260
rect 381 226 387 260
rect 341 201 387 226
rect 470 260 516 285
rect 470 226 476 260
rect 510 226 516 260
rect 470 201 516 226
rect 558 260 604 285
rect 558 226 564 260
rect 598 226 604 260
rect 558 201 604 226
rect 646 260 692 285
rect 646 226 652 260
rect 686 226 692 260
rect 646 201 692 226
rect 776 260 822 285
rect 776 226 782 260
rect 816 226 822 260
rect 776 201 822 226
rect 864 260 910 285
rect 864 226 870 260
rect 904 226 910 260
rect 864 201 910 226
rect 952 260 998 285
rect 952 226 958 260
rect 992 226 998 260
rect 952 201 998 226
rect 1040 260 1086 285
rect 1040 226 1046 260
rect 1080 226 1086 260
rect 1040 201 1086 226
rect 1128 260 1174 285
rect 1128 226 1134 260
rect 1168 226 1174 260
rect 1128 201 1174 226
rect 1216 260 1262 285
rect 1216 226 1222 260
rect 1256 226 1262 260
rect 1216 201 1262 226
rect 259 172 293 201
rect 476 172 510 201
rect 782 172 816 201
rect 958 172 992 201
rect 1134 172 1168 201
rect 99 138 1304 172
<< via1 >>
rect 99 1088 151 1140
rect 473 1053 525 1062
rect 473 1019 488 1053
rect 488 1019 522 1053
rect 522 1019 525 1053
rect 473 1010 525 1019
rect 1468 1106 1524 1162
rect 99 410 151 462
rect 473 357 525 366
rect 473 323 488 357
rect 488 323 522 357
rect 522 323 525 357
rect 473 314 525 323
rect 1562 410 1618 466
<< metal2 >>
rect 473 1391 526 1499
rect 99 1140 151 1150
rect 99 462 151 1088
rect 99 400 151 410
rect 473 1062 525 1391
rect 1468 1369 1524 1379
rect 1468 1162 1524 1313
rect 1468 1096 1524 1106
rect 1562 1243 1618 1253
rect 473 366 525 1010
rect 1562 466 1618 1187
rect 1562 376 1618 410
rect 473 0 525 314
<< via2 >>
rect 1468 1313 1524 1369
rect 1562 1187 1618 1243
<< metal3 >>
rect 1458 1369 2762 1374
rect 1458 1313 1468 1369
rect 1524 1313 2762 1369
rect 1458 1308 2762 1313
rect 1552 1243 2762 1248
rect 1552 1187 1562 1243
rect 1618 1187 2762 1243
rect 1552 1182 2762 1187
<< labels >>
rlabel metal1 0 1106 34 1140 0 A0
<< end >>
