magic
tech sky130A
magscale 1 2
timestamp 1702396496
<< error_p >>
rect -239 114 -181 120
rect 181 114 239 120
rect -239 80 -227 114
rect 181 80 193 114
rect -239 74 -181 80
rect 181 74 239 80
rect -449 -80 -391 -74
rect -29 -80 29 -74
rect 391 -80 449 -74
rect -449 -114 -437 -80
rect -29 -114 -17 -80
rect 391 -114 403 -80
rect -449 -120 -391 -114
rect -29 -120 29 -114
rect 391 -120 449 -114
<< nmos >>
rect -435 -42 -405 42
rect -225 -42 -195 42
rect -15 -42 15 42
rect 195 -42 225 42
rect 405 -42 435 42
<< ndiff >>
rect -497 30 -435 42
rect -497 -30 -485 30
rect -451 -30 -435 30
rect -497 -42 -435 -30
rect -405 30 -343 42
rect -405 -30 -389 30
rect -355 -30 -343 30
rect -405 -42 -343 -30
rect -287 30 -225 42
rect -287 -30 -275 30
rect -241 -30 -225 30
rect -287 -42 -225 -30
rect -195 30 -133 42
rect -195 -30 -179 30
rect -145 -30 -133 30
rect -195 -42 -133 -30
rect -77 30 -15 42
rect -77 -30 -65 30
rect -31 -30 -15 30
rect -77 -42 -15 -30
rect 15 30 77 42
rect 15 -30 31 30
rect 65 -30 77 30
rect 15 -42 77 -30
rect 133 30 195 42
rect 133 -30 145 30
rect 179 -30 195 30
rect 133 -42 195 -30
rect 225 30 287 42
rect 225 -30 241 30
rect 275 -30 287 30
rect 225 -42 287 -30
rect 343 30 405 42
rect 343 -30 355 30
rect 389 -30 405 30
rect 343 -42 405 -30
rect 435 30 497 42
rect 435 -30 451 30
rect 485 -30 497 30
rect 435 -42 497 -30
<< ndiffc >>
rect -485 -30 -451 30
rect -389 -30 -355 30
rect -275 -30 -241 30
rect -179 -30 -145 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 145 -30 179 30
rect 241 -30 275 30
rect 355 -30 389 30
rect 451 -30 485 30
<< poly >>
rect -243 114 -177 130
rect -243 80 -227 114
rect -193 80 -177 114
rect -435 42 -405 68
rect -243 64 -177 80
rect 177 114 243 130
rect 177 80 193 114
rect 227 80 243 114
rect -225 42 -195 64
rect -15 42 15 68
rect 177 64 243 80
rect 195 42 225 64
rect 405 42 435 68
rect -435 -64 -405 -42
rect -453 -80 -387 -64
rect -225 -68 -195 -42
rect -15 -64 15 -42
rect -453 -114 -437 -80
rect -403 -114 -387 -80
rect -453 -130 -387 -114
rect -33 -80 33 -64
rect 195 -68 225 -42
rect 405 -64 435 -42
rect -33 -114 -17 -80
rect 17 -114 33 -80
rect -33 -130 33 -114
rect 387 -80 453 -64
rect 387 -114 403 -80
rect 437 -114 453 -80
rect 387 -130 453 -114
<< polycont >>
rect -227 80 -193 114
rect 193 80 227 114
rect -437 -114 -403 -80
rect -17 -114 17 -80
rect 403 -114 437 -80
<< locali >>
rect -243 80 -227 114
rect -193 80 -177 114
rect 177 80 193 114
rect 227 80 243 114
rect -485 30 -451 46
rect -485 -46 -451 -30
rect -389 30 -355 46
rect -389 -46 -355 -30
rect -275 30 -241 46
rect -275 -46 -241 -30
rect -179 30 -145 46
rect -179 -46 -145 -30
rect -65 30 -31 46
rect -65 -46 -31 -30
rect 31 30 65 46
rect 31 -46 65 -30
rect 145 30 179 46
rect 145 -46 179 -30
rect 241 30 275 46
rect 241 -46 275 -30
rect 355 30 389 46
rect 355 -46 389 -30
rect 451 30 485 46
rect 451 -46 485 -30
rect -453 -114 -437 -80
rect -403 -114 -387 -80
rect -33 -114 -17 -80
rect 17 -114 33 -80
rect 387 -114 403 -80
rect 437 -114 453 -80
<< viali >>
rect -227 80 -193 114
rect 193 80 227 114
rect -485 -30 -451 30
rect -389 -30 -355 30
rect -275 -30 -241 30
rect -179 -30 -145 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 145 -30 179 30
rect 241 -30 275 30
rect 355 -30 389 30
rect 451 -30 485 30
rect -437 -114 -403 -80
rect -17 -114 17 -80
rect 403 -114 437 -80
<< metal1 >>
rect -239 114 -181 120
rect -239 80 -227 114
rect -193 80 -181 114
rect -239 74 -181 80
rect 181 114 239 120
rect 181 80 193 114
rect 227 80 239 114
rect 181 74 239 80
rect -491 30 -445 42
rect -491 -30 -485 30
rect -451 -30 -445 30
rect -491 -42 -445 -30
rect -395 30 -349 42
rect -395 -30 -389 30
rect -355 -30 -349 30
rect -395 -42 -349 -30
rect -281 30 -235 42
rect -281 -30 -275 30
rect -241 -30 -235 30
rect -281 -42 -235 -30
rect -185 30 -139 42
rect -185 -30 -179 30
rect -145 -30 -139 30
rect -185 -42 -139 -30
rect -71 30 -25 42
rect -71 -30 -65 30
rect -31 -30 -25 30
rect -71 -42 -25 -30
rect 25 30 71 42
rect 25 -30 31 30
rect 65 -30 71 30
rect 25 -42 71 -30
rect 139 30 185 42
rect 139 -30 145 30
rect 179 -30 185 30
rect 139 -42 185 -30
rect 235 30 281 42
rect 235 -30 241 30
rect 275 -30 281 30
rect 235 -42 281 -30
rect 349 30 395 42
rect 349 -30 355 30
rect 389 -30 395 30
rect 349 -42 395 -30
rect 445 30 491 42
rect 445 -30 451 30
rect 485 -30 491 30
rect 445 -42 491 -30
rect -449 -80 -391 -74
rect -449 -114 -437 -80
rect -403 -114 -391 -80
rect -449 -120 -391 -114
rect -29 -80 29 -74
rect -29 -114 -17 -80
rect 17 -114 29 -80
rect -29 -120 29 -114
rect 391 -80 449 -74
rect 391 -114 403 -80
rect 437 -114 449 -80
rect 391 -120 449 -114
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 5 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
