magic
tech sky130A
magscale 1 2
timestamp 1702727116
<< nwell >>
rect 338 1619 644 1848
rect 0 1116 720 1619
rect 187 337 545 661
<< nmos >>
rect 94 2034 124 2202
rect 432 1954 462 2354
rect 520 1954 550 2354
rect 94 1688 124 1772
rect 182 1688 212 1772
rect 93 828 123 948
rect 293 828 323 988
rect 381 828 411 988
rect 595 828 625 948
rect 421 69 451 269
<< pmos >>
rect 94 1473 124 1557
rect 182 1473 212 1557
rect 432 1386 462 1786
rect 520 1386 550 1786
rect 293 1178 323 1262
rect 381 1178 411 1262
rect 421 399 451 599
<< ndiff >>
rect 374 2342 432 2354
rect 36 2190 94 2202
rect 36 2046 48 2190
rect 82 2046 94 2190
rect 36 2034 94 2046
rect 124 2190 182 2202
rect 124 2046 136 2190
rect 170 2046 182 2190
rect 124 2034 182 2046
rect 374 1966 386 2342
rect 420 1966 432 2342
rect 374 1954 432 1966
rect 462 2342 520 2354
rect 462 1966 474 2342
rect 508 1966 520 2342
rect 462 1954 520 1966
rect 550 2342 608 2354
rect 550 1966 562 2342
rect 596 1966 608 2342
rect 550 1954 608 1966
rect 36 1760 94 1772
rect 36 1700 48 1760
rect 82 1700 94 1760
rect 36 1688 94 1700
rect 124 1760 182 1772
rect 124 1700 136 1760
rect 170 1700 182 1760
rect 124 1688 182 1700
rect 212 1760 270 1772
rect 212 1700 224 1760
rect 258 1700 270 1760
rect 212 1688 270 1700
rect 235 976 293 988
rect 35 936 93 948
rect 35 840 47 936
rect 81 840 93 936
rect 35 828 93 840
rect 123 936 181 948
rect 123 840 135 936
rect 169 840 181 936
rect 123 828 181 840
rect 235 840 247 976
rect 281 840 293 976
rect 235 828 293 840
rect 323 976 381 988
rect 323 840 335 976
rect 369 840 381 976
rect 323 828 381 840
rect 411 976 469 988
rect 411 840 423 976
rect 457 840 469 976
rect 411 828 469 840
rect 537 936 595 948
rect 537 840 549 936
rect 583 840 595 936
rect 537 828 595 840
rect 625 936 683 948
rect 625 840 637 936
rect 671 840 683 936
rect 625 828 683 840
rect 363 257 421 269
rect 363 81 375 257
rect 409 81 421 257
rect 363 69 421 81
rect 451 257 509 269
rect 451 81 463 257
rect 497 81 509 257
rect 451 69 509 81
<< pdiff >>
rect 374 1774 432 1786
rect 36 1545 94 1557
rect 36 1485 48 1545
rect 82 1485 94 1545
rect 36 1473 94 1485
rect 124 1545 182 1557
rect 124 1485 136 1545
rect 170 1485 182 1545
rect 124 1473 182 1485
rect 212 1545 270 1557
rect 212 1485 224 1545
rect 258 1485 270 1545
rect 212 1473 270 1485
rect 374 1398 386 1774
rect 420 1398 432 1774
rect 374 1386 432 1398
rect 462 1774 520 1786
rect 462 1398 474 1774
rect 508 1398 520 1774
rect 462 1386 520 1398
rect 550 1774 608 1786
rect 550 1398 562 1774
rect 596 1398 608 1774
rect 550 1386 608 1398
rect 235 1250 293 1262
rect 235 1190 247 1250
rect 281 1190 293 1250
rect 235 1178 293 1190
rect 323 1250 381 1262
rect 323 1190 335 1250
rect 369 1190 381 1250
rect 323 1178 381 1190
rect 411 1250 469 1262
rect 411 1190 423 1250
rect 457 1190 469 1250
rect 411 1178 469 1190
rect 363 587 421 599
rect 363 411 375 587
rect 409 411 421 587
rect 363 399 421 411
rect 451 587 509 599
rect 451 411 463 587
rect 497 411 509 587
rect 451 399 509 411
<< ndiffc >>
rect 48 2046 82 2190
rect 136 2046 170 2190
rect 386 1966 420 2342
rect 474 1966 508 2342
rect 562 1966 596 2342
rect 48 1700 82 1760
rect 136 1700 170 1760
rect 224 1700 258 1760
rect 47 840 81 936
rect 135 840 169 936
rect 247 840 281 976
rect 335 840 369 976
rect 423 840 457 976
rect 549 840 583 936
rect 637 840 671 936
rect 375 81 409 257
rect 463 81 497 257
<< pdiffc >>
rect 48 1485 82 1545
rect 136 1485 170 1545
rect 224 1485 258 1545
rect 386 1398 420 1774
rect 474 1398 508 1774
rect 562 1398 596 1774
rect 247 1190 281 1250
rect 335 1190 369 1250
rect 423 1190 457 1250
rect 375 411 409 587
rect 463 411 497 587
<< psubdiff >>
rect 237 2329 319 2353
rect 237 2295 262 2329
rect 296 2295 319 2329
rect 237 2271 319 2295
rect 310 750 392 774
rect 310 716 335 750
rect 369 716 392 750
rect 310 692 392 716
<< nsubdiff >>
rect 523 1250 605 1262
rect 523 1190 547 1250
rect 581 1190 605 1250
rect 523 1178 605 1190
rect 223 523 305 535
rect 223 463 247 523
rect 281 463 305 523
rect 223 451 305 463
<< psubdiffcont >>
rect 262 2295 296 2329
rect 335 716 369 750
<< nsubdiffcont >>
rect 547 1190 581 1250
rect 247 463 281 523
<< poly >>
rect 432 2354 462 2380
rect 520 2354 550 2380
rect 94 2305 193 2321
rect 94 2271 143 2305
rect 177 2271 193 2305
rect 94 2255 193 2271
rect 94 2228 125 2255
rect 94 2202 124 2228
rect 94 2008 124 2034
rect 262 1996 328 2007
rect 262 1982 278 1996
rect 182 1962 278 1982
rect 312 1962 328 1996
rect 182 1952 328 1962
rect 39 1909 124 1925
rect 39 1875 55 1909
rect 89 1875 124 1909
rect 39 1859 124 1875
rect 94 1772 124 1859
rect 182 1772 212 1952
rect 286 1882 352 1898
rect 432 1882 462 1954
rect 286 1848 302 1882
rect 336 1848 462 1882
rect 286 1832 352 1848
rect 432 1786 462 1848
rect 520 1923 550 1954
rect 520 1907 600 1923
rect 520 1873 550 1907
rect 584 1873 600 1907
rect 520 1858 600 1873
rect 520 1786 550 1858
rect 94 1662 124 1688
rect 182 1662 212 1688
rect 94 1557 124 1583
rect 182 1557 212 1583
rect 94 1447 124 1473
rect 182 1447 212 1473
rect 94 1411 212 1447
rect 120 1377 136 1411
rect 170 1377 186 1411
rect 120 1361 186 1377
rect 432 1360 462 1386
rect 520 1360 550 1386
rect 293 1262 323 1288
rect 381 1262 411 1288
rect 293 1143 323 1178
rect 257 1131 323 1143
rect 257 1097 273 1131
rect 307 1097 323 1131
rect 257 1086 323 1097
rect 27 1063 123 1079
rect 27 1029 43 1063
rect 77 1029 123 1063
rect 27 1013 123 1029
rect 93 948 123 1013
rect 293 988 323 1086
rect 381 1075 411 1178
rect 381 1060 447 1075
rect 381 1026 397 1060
rect 431 1026 447 1060
rect 381 1009 447 1026
rect 578 1063 644 1079
rect 578 1029 594 1063
rect 628 1029 644 1063
rect 578 1013 644 1029
rect 381 988 411 1009
rect 595 948 625 1013
rect 93 802 123 828
rect 293 802 323 828
rect 381 802 411 828
rect 595 802 625 828
rect 421 599 451 625
rect 421 352 451 399
rect 538 352 593 368
rect 421 318 549 352
rect 583 318 593 352
rect 421 269 451 318
rect 538 302 593 318
rect 421 43 451 69
<< polycont >>
rect 143 2271 177 2305
rect 278 1962 312 1996
rect 55 1875 89 1909
rect 302 1848 336 1882
rect 550 1873 584 1907
rect 136 1377 170 1411
rect 273 1097 307 1131
rect 43 1029 77 1063
rect 397 1026 431 1060
rect 594 1029 628 1063
rect 549 318 583 352
<< locali >>
rect 143 2305 177 2488
rect 237 2329 319 2353
rect 237 2295 262 2329
rect 296 2295 319 2329
rect 237 2271 319 2295
rect 386 2342 420 2358
rect 143 2255 177 2271
rect 48 2190 82 2206
rect 48 2030 82 2046
rect 136 2190 170 2206
rect 136 2030 170 2046
rect 262 1962 278 1996
rect 312 1962 328 1996
rect 39 1875 55 1909
rect 89 1875 105 1909
rect 386 1907 420 1966
rect 474 2342 508 2358
rect 474 1950 508 1966
rect 562 2342 596 2358
rect 596 1966 668 1984
rect 562 1950 668 1966
rect 224 1848 302 1882
rect 336 1848 352 1882
rect 386 1873 550 1907
rect 584 1873 600 1907
rect 48 1760 82 1776
rect 48 1545 82 1700
rect 136 1760 170 1776
rect 136 1684 170 1700
rect 224 1760 258 1848
rect 48 1411 82 1485
rect 136 1545 170 1561
rect 136 1469 170 1485
rect 224 1545 258 1700
rect 224 1469 258 1485
rect 386 1774 420 1873
rect 634 1791 668 1950
rect 48 1377 136 1411
rect 170 1377 186 1411
rect 386 1338 420 1398
rect 474 1774 508 1790
rect 474 1382 508 1398
rect 562 1774 668 1791
rect 596 1757 668 1774
rect 562 1382 596 1398
rect 46 1304 420 1338
rect 46 1227 80 1304
rect 247 1250 281 1266
rect 189 1190 247 1208
rect 189 1174 281 1190
rect 335 1250 369 1266
rect 335 1174 369 1190
rect 423 1250 457 1266
rect 27 1029 34 1063
rect 86 1029 93 1063
rect 189 1060 223 1174
rect 423 1131 457 1190
rect 547 1250 581 1274
rect 547 1166 581 1190
rect 257 1097 273 1131
rect 307 1097 515 1131
rect 135 1026 397 1060
rect 431 1026 447 1060
rect 47 936 81 952
rect 47 824 81 840
rect 135 936 169 1026
rect 135 824 169 840
rect 247 976 281 1026
rect 481 992 515 1097
rect 578 1029 585 1063
rect 637 1029 644 1063
rect 247 824 281 840
rect 335 976 369 992
rect 335 824 369 840
rect 423 976 583 992
rect 457 958 583 976
rect 423 824 457 840
rect 549 936 583 958
rect 310 750 392 774
rect 310 716 335 750
rect 369 716 392 750
rect 310 692 392 716
rect 375 587 409 603
rect 247 523 281 547
rect 281 477 375 511
rect 247 439 281 463
rect 375 395 409 411
rect 463 587 497 603
rect 463 395 497 411
rect 549 352 583 840
rect 637 936 671 952
rect 637 824 671 840
rect 549 297 583 318
rect 375 257 409 273
rect 375 65 409 81
rect 463 257 497 273
rect 463 65 497 81
<< viali >>
rect 143 2488 177 2522
rect 262 2295 296 2329
rect 48 2046 82 2190
rect 136 2046 170 2190
rect 278 1962 312 1996
rect 386 1966 420 2342
rect 55 1875 89 1909
rect 474 1966 508 2342
rect 562 1966 596 2342
rect 48 1700 82 1760
rect 136 1700 170 1760
rect 224 1700 258 1760
rect 48 1485 82 1545
rect 136 1485 170 1545
rect 224 1485 258 1545
rect 386 1398 420 1774
rect 474 1398 508 1774
rect 562 1398 596 1774
rect 46 1193 80 1227
rect 247 1190 281 1250
rect 335 1190 369 1250
rect 423 1190 457 1250
rect 34 1063 86 1081
rect 34 1029 43 1063
rect 43 1029 77 1063
rect 77 1029 86 1063
rect 547 1190 581 1250
rect 47 840 81 936
rect 135 840 169 936
rect 585 1063 637 1081
rect 585 1029 594 1063
rect 594 1029 628 1063
rect 628 1029 637 1063
rect 247 840 281 976
rect 335 840 369 976
rect 423 840 457 976
rect 549 840 583 936
rect 335 716 369 750
rect 375 411 409 587
rect 463 411 497 587
rect 637 840 671 936
rect 375 81 409 257
rect 463 81 497 257
<< metal1 >>
rect 316 2614 326 2632
rect 0 2580 326 2614
rect 378 2614 388 2632
rect 378 2580 720 2614
rect 131 2522 189 2528
rect 234 2522 244 2540
rect 0 2488 143 2522
rect 177 2488 244 2522
rect 296 2522 306 2540
rect 296 2488 720 2522
rect 131 2482 189 2488
rect 396 2427 406 2445
rect 0 2393 406 2427
rect 458 2427 468 2445
rect 458 2393 720 2427
rect 48 2202 82 2393
rect 237 2329 309 2393
rect 474 2354 508 2393
rect 237 2295 262 2329
rect 296 2295 309 2329
rect 237 2271 309 2295
rect 380 2342 426 2354
rect 42 2190 88 2202
rect 42 2046 48 2190
rect 82 2046 88 2190
rect 42 2034 88 2046
rect 130 2190 176 2202
rect 130 2046 136 2190
rect 170 2046 176 2190
rect 130 2034 176 2046
rect 36 1866 46 1918
rect 98 1866 108 1918
rect 136 1772 170 2034
rect 266 1996 324 2002
rect 266 1962 278 1996
rect 312 1962 324 1996
rect 266 1956 324 1962
rect 380 1966 386 2342
rect 420 1966 426 2342
rect 278 1901 312 1956
rect 380 1954 426 1966
rect 468 2342 514 2354
rect 468 1966 474 2342
rect 508 1966 514 2342
rect 468 1954 514 1966
rect 556 2342 602 2354
rect 556 1966 562 2342
rect 596 1966 602 2342
rect 556 1954 602 1966
rect 630 1901 640 1910
rect 278 1867 640 1901
rect 630 1858 640 1867
rect 692 1858 702 1910
rect 380 1774 426 1786
rect 42 1760 88 1772
rect 42 1700 48 1760
rect 82 1700 88 1760
rect 42 1688 88 1700
rect 130 1760 176 1772
rect 130 1700 136 1760
rect 170 1700 176 1760
rect 130 1688 176 1700
rect 218 1760 264 1772
rect 218 1700 224 1760
rect 258 1700 264 1760
rect 218 1688 264 1700
rect 42 1545 88 1557
rect 42 1485 48 1545
rect 82 1485 88 1545
rect 42 1473 88 1485
rect 130 1545 176 1557
rect 130 1485 136 1545
rect 170 1485 176 1545
rect 130 1473 176 1485
rect 218 1545 264 1557
rect 218 1485 224 1545
rect 258 1485 264 1545
rect 218 1473 264 1485
rect 135 1324 170 1473
rect 380 1398 386 1774
rect 420 1398 426 1774
rect 380 1386 426 1398
rect 468 1774 514 1786
rect 468 1398 474 1774
rect 508 1398 514 1774
rect 468 1386 514 1398
rect 556 1774 602 1786
rect 556 1398 562 1774
rect 596 1439 602 1774
rect 596 1398 628 1439
rect 556 1387 628 1398
rect 680 1387 690 1439
rect 556 1386 690 1387
rect 316 1324 326 1342
rect 0 1290 326 1324
rect 378 1324 388 1342
rect 474 1324 509 1386
rect 378 1290 720 1324
rect 335 1262 369 1290
rect 547 1262 581 1290
rect 241 1250 287 1262
rect 27 1184 37 1236
rect 90 1184 100 1236
rect 241 1190 247 1250
rect 281 1190 287 1250
rect 241 1178 287 1190
rect 329 1250 375 1262
rect 329 1190 335 1250
rect 369 1190 375 1250
rect 329 1178 375 1190
rect 417 1250 463 1262
rect 417 1190 423 1250
rect 457 1190 463 1250
rect 417 1178 463 1190
rect 541 1250 587 1262
rect 541 1190 547 1250
rect 581 1190 587 1250
rect 541 1178 587 1190
rect 22 1081 98 1087
rect 22 1029 34 1081
rect 86 1072 98 1081
rect 234 1072 244 1090
rect 86 1038 244 1072
rect 296 1072 306 1090
rect 573 1081 649 1087
rect 573 1072 585 1081
rect 296 1038 585 1072
rect 86 1029 98 1038
rect 22 1023 98 1029
rect 573 1029 585 1038
rect 637 1029 649 1081
rect 573 1023 649 1029
rect 241 976 287 988
rect 41 936 87 948
rect 41 886 47 936
rect 81 886 87 936
rect 129 936 175 948
rect 28 834 38 886
rect 90 834 100 886
rect 129 840 135 936
rect 169 840 175 936
rect 41 828 87 834
rect 129 828 175 840
rect 241 840 247 976
rect 281 840 287 976
rect 241 828 287 840
rect 329 976 375 988
rect 329 840 335 976
rect 369 840 375 976
rect 329 828 375 840
rect 417 976 463 988
rect 417 840 423 976
rect 457 840 463 976
rect 417 828 463 840
rect 543 936 589 948
rect 543 840 549 936
rect 583 840 589 936
rect 631 936 677 948
rect 631 886 637 936
rect 671 886 677 936
rect 543 828 589 840
rect 618 834 628 886
rect 680 834 690 886
rect 631 828 677 834
rect 335 800 369 828
rect 0 766 406 800
rect 249 269 283 766
rect 323 750 406 766
rect 323 716 335 750
rect 369 748 406 750
rect 458 766 720 800
rect 458 748 468 766
rect 369 716 382 748
rect 323 711 382 716
rect 323 710 381 711
rect 316 616 326 669
rect 378 616 415 669
rect 316 599 415 616
rect 369 587 415 599
rect 369 411 375 587
rect 409 411 415 587
rect 369 399 415 411
rect 457 587 503 599
rect 457 411 463 587
rect 497 411 503 587
rect 457 399 503 411
rect 463 269 497 399
rect 249 257 415 269
rect 249 235 375 257
rect 369 81 375 235
rect 409 81 415 257
rect 369 69 415 81
rect 457 257 503 269
rect 457 81 463 257
rect 497 81 503 257
rect 457 69 503 81
rect 463 0 497 69
<< via1 >>
rect 326 2580 378 2632
rect 244 2488 296 2540
rect 406 2393 458 2445
rect 46 1909 98 1918
rect 46 1875 55 1909
rect 55 1875 89 1909
rect 89 1875 98 1909
rect 46 1866 98 1875
rect 640 1858 692 1910
rect 628 1387 680 1439
rect 326 1290 378 1342
rect 37 1227 90 1236
rect 37 1193 46 1227
rect 46 1193 80 1227
rect 80 1193 90 1227
rect 37 1184 90 1193
rect 244 1038 296 1090
rect 38 840 47 886
rect 47 840 81 886
rect 81 840 90 886
rect 38 834 90 840
rect 628 840 637 886
rect 637 840 671 886
rect 671 840 680 886
rect 628 834 680 840
rect 406 748 458 800
rect 326 616 378 669
<< metal2 >>
rect 12 2468 64 2666
rect 12 2434 98 2468
rect 46 1918 98 2434
rect 46 1856 98 1866
rect 38 1246 90 1324
rect 37 1236 90 1246
rect 37 1174 90 1184
rect 38 886 90 1174
rect 38 828 90 834
rect 164 0 216 2666
rect 326 2632 378 2639
rect 244 2540 296 2550
rect 244 1090 296 2488
rect 244 1028 296 1038
rect 326 1342 378 2580
rect 326 669 378 1290
rect 406 2445 458 2455
rect 406 800 458 2393
rect 406 738 458 748
rect 326 606 378 616
rect 488 0 540 2667
rect 640 1910 692 2666
rect 640 1848 692 1858
rect 628 1439 680 1449
rect 628 886 680 1387
rect 628 828 680 834
<< labels >>
rlabel metal2 12 2614 64 2666 0 DR_
rlabel metal2 164 2614 216 2666 0 DW_
rlabel metal2 488 2615 540 2667 0 DW
rlabel metal2 640 2614 692 2666 0 DR
rlabel metal1 12 2580 46 2614 0 VDD
rlabel metal1 12 2488 46 2522 0 SAEN
rlabel metal1 12 2393 46 2427 0 VSS
rlabel metal2 164 0 216 52 0 DW_
rlabel metal2 488 0 540 52 0 DW
rlabel metal1 463 0 497 34 0 SB
rlabel metal1 0 1290 34 1324 0 VDD
rlabel metal1 0 766 34 800 0 VSS
<< end >>
