magic
tech sky130A
magscale 1 2
timestamp 1702831315
<< nwell >>
rect 2806 1876 3136 1877
rect 0 1669 3136 1876
rect 0 1668 2806 1669
rect 0 1214 3242 1290
rect 0 1082 3460 1214
rect 2806 1006 3460 1082
rect 0 350 3719 558
rect 1420 137 1638 350
<< pwell >>
rect 10 1491 120 1503
rect 2486 1491 2596 1503
rect 2816 1492 2926 1504
rect 10 1355 320 1491
rect 2180 1355 2466 1491
rect 2486 1355 2796 1491
rect 2816 1356 3126 1492
rect 10 1343 120 1355
rect 2486 1343 2596 1355
rect 2816 1344 2926 1356
rect 2486 905 2596 917
rect 2180 769 2466 905
rect 2486 769 2796 905
rect 2486 757 2596 769
rect 338 173 448 185
rect 338 37 648 173
rect 808 37 1094 173
rect 1745 173 1855 185
rect 2612 173 2722 185
rect 3399 173 3509 185
rect 1745 37 2055 173
rect 2218 37 2592 173
rect 2612 37 2922 173
rect 3093 37 3379 173
rect 3399 37 3709 173
rect 338 25 448 37
rect 1745 25 1855 37
rect 2612 25 2722 37
rect 3399 25 3509 37
<< nmos >>
rect 206 1381 236 1465
rect 517 1381 547 1465
rect 605 1381 635 1465
rect 823 1381 853 1465
rect 911 1381 941 1465
rect 1129 1381 1159 1465
rect 1217 1381 1247 1465
rect 1434 1381 1465 1465
rect 1522 1381 1552 1465
rect 1740 1381 1770 1465
rect 1828 1381 1858 1465
rect 2046 1381 2076 1465
rect 2264 1381 2294 1465
rect 2352 1381 2382 1465
rect 2682 1381 2712 1465
rect 3012 1382 3042 1466
rect 517 795 547 879
rect 605 795 635 879
rect 823 795 853 879
rect 911 795 941 879
rect 1129 795 1159 879
rect 1217 795 1247 879
rect 1434 795 1465 879
rect 1522 795 1552 879
rect 1740 795 1770 879
rect 1828 795 1858 879
rect 2046 795 2076 879
rect 2264 795 2294 879
rect 2352 795 2382 879
rect 2682 795 2712 879
rect 2900 694 2930 854
rect 3118 694 3148 854
rect 3336 770 3366 854
rect 3547 694 3577 854
rect 534 63 564 147
rect 892 63 922 147
rect 980 63 1010 147
rect 1941 63 1971 147
rect 2302 63 2332 147
rect 2390 63 2420 147
rect 2478 63 2508 147
rect 2808 63 2838 147
rect 3177 63 3207 147
rect 3265 63 3295 147
rect 3595 63 3625 147
<< pmos >>
rect 206 1730 236 1814
rect 517 1730 547 1814
rect 605 1730 635 1814
rect 823 1730 853 1814
rect 911 1730 941 1814
rect 1129 1730 1159 1814
rect 1217 1730 1247 1814
rect 1434 1730 1465 1814
rect 1522 1730 1552 1814
rect 1740 1730 1770 1814
rect 1828 1730 1858 1814
rect 2046 1730 2076 1814
rect 2264 1730 2294 1814
rect 2352 1730 2382 1814
rect 2682 1730 2712 1814
rect 3012 1731 3042 1815
rect 517 1144 547 1228
rect 605 1144 635 1228
rect 823 1144 853 1228
rect 911 1144 941 1228
rect 1129 1144 1159 1228
rect 1217 1144 1247 1228
rect 1434 1144 1465 1228
rect 1522 1144 1552 1228
rect 1740 1144 1770 1228
rect 1828 1144 1858 1228
rect 2046 1144 2076 1228
rect 2264 1144 2294 1228
rect 2352 1144 2382 1228
rect 2682 1144 2712 1228
rect 2900 1068 2930 1228
rect 3118 1068 3148 1228
rect 3336 1068 3366 1152
rect 534 412 564 496
rect 892 412 922 496
rect 980 412 1010 496
rect 1470 412 1500 496
rect 1558 412 1588 496
rect 1941 412 1971 496
rect 2302 412 2332 496
rect 2390 412 2420 496
rect 2478 412 2508 496
rect 1514 199 1544 283
rect 2808 412 2838 496
rect 3177 412 3207 496
rect 3265 412 3295 496
rect 3595 412 3625 496
<< ndiff >>
rect 148 1440 206 1465
rect 148 1406 160 1440
rect 194 1406 206 1440
rect 148 1381 206 1406
rect 236 1440 294 1465
rect 236 1406 248 1440
rect 282 1406 294 1440
rect 236 1381 294 1406
rect 459 1453 517 1465
rect 459 1393 471 1453
rect 505 1393 517 1453
rect 459 1381 517 1393
rect 547 1453 605 1465
rect 547 1393 559 1453
rect 593 1393 605 1453
rect 547 1381 605 1393
rect 635 1453 693 1465
rect 635 1393 647 1453
rect 681 1393 693 1453
rect 635 1381 693 1393
rect 765 1453 823 1465
rect 765 1393 777 1453
rect 811 1393 823 1453
rect 765 1381 823 1393
rect 853 1453 911 1465
rect 853 1393 865 1453
rect 899 1393 911 1453
rect 853 1381 911 1393
rect 941 1453 999 1465
rect 941 1393 953 1453
rect 987 1393 999 1453
rect 941 1381 999 1393
rect 1071 1453 1129 1465
rect 1071 1393 1083 1453
rect 1117 1393 1129 1453
rect 1071 1381 1129 1393
rect 1159 1453 1217 1465
rect 1159 1393 1171 1453
rect 1205 1393 1217 1453
rect 1159 1381 1217 1393
rect 1247 1453 1305 1465
rect 1247 1393 1259 1453
rect 1293 1393 1305 1453
rect 1247 1381 1305 1393
rect 1376 1453 1434 1465
rect 1376 1393 1388 1453
rect 1422 1393 1434 1453
rect 1376 1381 1434 1393
rect 1465 1453 1522 1465
rect 1465 1393 1476 1453
rect 1510 1393 1522 1453
rect 1465 1381 1522 1393
rect 1552 1453 1610 1465
rect 1552 1393 1564 1453
rect 1598 1393 1610 1453
rect 1552 1381 1610 1393
rect 1682 1453 1740 1465
rect 1682 1393 1694 1453
rect 1728 1393 1740 1453
rect 1682 1381 1740 1393
rect 1770 1453 1828 1465
rect 1770 1393 1782 1453
rect 1816 1393 1828 1453
rect 1770 1381 1828 1393
rect 1858 1453 1916 1465
rect 1858 1393 1870 1453
rect 1904 1393 1916 1453
rect 1858 1381 1916 1393
rect 1988 1453 2046 1465
rect 1988 1393 2000 1453
rect 2034 1393 2046 1453
rect 1988 1381 2046 1393
rect 2076 1453 2134 1465
rect 2076 1393 2088 1453
rect 2122 1393 2134 1453
rect 2076 1381 2134 1393
rect 2206 1440 2264 1465
rect 2206 1406 2218 1440
rect 2252 1406 2264 1440
rect 2206 1381 2264 1406
rect 2294 1440 2352 1465
rect 2294 1406 2306 1440
rect 2340 1406 2352 1440
rect 2294 1381 2352 1406
rect 2382 1440 2440 1465
rect 2382 1406 2394 1440
rect 2428 1406 2440 1440
rect 2382 1381 2440 1406
rect 2624 1440 2682 1465
rect 2624 1406 2636 1440
rect 2670 1406 2682 1440
rect 2624 1381 2682 1406
rect 2712 1440 2770 1465
rect 2712 1406 2724 1440
rect 2758 1406 2770 1440
rect 2712 1381 2770 1406
rect 2954 1441 3012 1466
rect 2954 1407 2966 1441
rect 3000 1407 3012 1441
rect 2954 1382 3012 1407
rect 3042 1441 3100 1466
rect 3042 1407 3054 1441
rect 3088 1407 3100 1441
rect 3042 1382 3100 1407
rect 459 867 517 879
rect 459 807 471 867
rect 505 807 517 867
rect 459 795 517 807
rect 547 867 605 879
rect 547 807 559 867
rect 593 807 605 867
rect 547 795 605 807
rect 635 867 693 879
rect 635 807 647 867
rect 681 807 693 867
rect 635 795 693 807
rect 765 867 823 879
rect 765 807 777 867
rect 811 807 823 867
rect 765 795 823 807
rect 853 867 911 879
rect 853 807 865 867
rect 899 807 911 867
rect 853 795 911 807
rect 941 867 999 879
rect 941 807 953 867
rect 987 807 999 867
rect 941 795 999 807
rect 1071 867 1129 879
rect 1071 807 1083 867
rect 1117 807 1129 867
rect 1071 795 1129 807
rect 1159 867 1217 879
rect 1159 807 1171 867
rect 1205 807 1217 867
rect 1159 795 1217 807
rect 1247 867 1305 879
rect 1247 807 1259 867
rect 1293 807 1305 867
rect 1247 795 1305 807
rect 1376 867 1434 879
rect 1376 807 1388 867
rect 1422 807 1434 867
rect 1376 795 1434 807
rect 1465 867 1522 879
rect 1465 807 1476 867
rect 1510 807 1522 867
rect 1465 795 1522 807
rect 1552 867 1610 879
rect 1552 807 1564 867
rect 1598 807 1610 867
rect 1552 795 1610 807
rect 1682 867 1740 879
rect 1682 807 1694 867
rect 1728 807 1740 867
rect 1682 795 1740 807
rect 1770 867 1828 879
rect 1770 807 1782 867
rect 1816 807 1828 867
rect 1770 795 1828 807
rect 1858 867 1916 879
rect 1858 807 1870 867
rect 1904 807 1916 867
rect 1858 795 1916 807
rect 1988 867 2046 879
rect 1988 807 2000 867
rect 2034 807 2046 867
rect 1988 795 2046 807
rect 2076 867 2134 879
rect 2076 807 2088 867
rect 2122 807 2134 867
rect 2076 795 2134 807
rect 2206 854 2264 879
rect 2206 820 2218 854
rect 2252 820 2264 854
rect 2206 795 2264 820
rect 2294 854 2352 879
rect 2294 820 2306 854
rect 2340 820 2352 854
rect 2294 795 2352 820
rect 2382 854 2440 879
rect 2382 820 2394 854
rect 2428 820 2440 854
rect 2382 795 2440 820
rect 2624 854 2682 879
rect 2624 820 2636 854
rect 2670 820 2682 854
rect 2624 795 2682 820
rect 2712 854 2770 879
rect 2712 820 2724 854
rect 2758 820 2770 854
rect 2712 795 2770 820
rect 2842 842 2900 854
rect 2842 706 2854 842
rect 2888 706 2900 842
rect 2842 694 2900 706
rect 2930 842 2988 854
rect 2930 706 2942 842
rect 2976 706 2988 842
rect 2930 694 2988 706
rect 3060 842 3118 854
rect 3060 706 3072 842
rect 3106 706 3118 842
rect 3060 694 3118 706
rect 3148 842 3206 854
rect 3148 706 3160 842
rect 3194 706 3206 842
rect 3278 842 3336 854
rect 3278 782 3290 842
rect 3324 782 3336 842
rect 3278 770 3336 782
rect 3366 842 3424 854
rect 3366 782 3378 842
rect 3412 782 3424 842
rect 3366 770 3424 782
rect 3489 842 3547 854
rect 3148 694 3206 706
rect 3489 706 3501 842
rect 3535 706 3547 842
rect 3489 694 3547 706
rect 3577 842 3635 854
rect 3577 706 3589 842
rect 3623 706 3635 842
rect 3577 694 3635 706
rect 476 122 534 147
rect 476 88 488 122
rect 522 88 534 122
rect 476 63 534 88
rect 564 122 622 147
rect 564 88 576 122
rect 610 88 622 122
rect 564 63 622 88
rect 834 122 892 147
rect 834 88 846 122
rect 880 88 892 122
rect 834 63 892 88
rect 922 122 980 147
rect 922 88 934 122
rect 968 88 980 122
rect 922 63 980 88
rect 1010 122 1068 147
rect 1010 88 1022 122
rect 1056 88 1068 122
rect 1010 63 1068 88
rect 1883 122 1941 147
rect 1883 88 1895 122
rect 1929 88 1941 122
rect 1883 63 1941 88
rect 1971 122 2029 147
rect 1971 88 1983 122
rect 2017 88 2029 122
rect 1971 63 2029 88
rect 2244 122 2302 147
rect 2244 88 2256 122
rect 2290 88 2302 122
rect 2244 63 2302 88
rect 2332 122 2390 147
rect 2332 88 2344 122
rect 2378 88 2390 122
rect 2332 63 2390 88
rect 2420 122 2478 147
rect 2420 88 2432 122
rect 2466 88 2478 122
rect 2420 63 2478 88
rect 2508 122 2566 147
rect 2508 88 2520 122
rect 2554 88 2566 122
rect 2508 63 2566 88
rect 2750 122 2808 147
rect 2750 88 2762 122
rect 2796 88 2808 122
rect 2750 63 2808 88
rect 2838 122 2896 147
rect 2838 88 2850 122
rect 2884 88 2896 122
rect 2838 63 2896 88
rect 3119 122 3177 147
rect 3119 88 3131 122
rect 3165 88 3177 122
rect 3119 63 3177 88
rect 3207 122 3265 147
rect 3207 88 3219 122
rect 3253 88 3265 122
rect 3207 63 3265 88
rect 3295 122 3353 147
rect 3295 88 3307 122
rect 3341 88 3353 122
rect 3295 63 3353 88
rect 3537 122 3595 147
rect 3537 88 3549 122
rect 3583 88 3595 122
rect 3537 63 3595 88
rect 3625 122 3683 147
rect 3625 88 3637 122
rect 3671 88 3683 122
rect 3625 63 3683 88
<< pdiff >>
rect 148 1789 206 1814
rect 148 1755 160 1789
rect 194 1755 206 1789
rect 148 1730 206 1755
rect 236 1789 294 1814
rect 236 1755 248 1789
rect 282 1755 294 1789
rect 236 1730 294 1755
rect 459 1802 517 1814
rect 459 1742 471 1802
rect 505 1742 517 1802
rect 459 1730 517 1742
rect 547 1802 605 1814
rect 547 1742 559 1802
rect 593 1742 605 1802
rect 547 1730 605 1742
rect 635 1802 693 1814
rect 635 1742 647 1802
rect 681 1742 693 1802
rect 635 1730 693 1742
rect 765 1802 823 1814
rect 765 1742 777 1802
rect 811 1742 823 1802
rect 765 1730 823 1742
rect 853 1802 911 1814
rect 853 1742 865 1802
rect 899 1742 911 1802
rect 853 1730 911 1742
rect 941 1802 999 1814
rect 941 1742 953 1802
rect 987 1742 999 1802
rect 941 1730 999 1742
rect 1071 1802 1129 1814
rect 1071 1742 1083 1802
rect 1117 1742 1129 1802
rect 1071 1730 1129 1742
rect 1159 1802 1217 1814
rect 1159 1742 1171 1802
rect 1205 1742 1217 1802
rect 1159 1730 1217 1742
rect 1247 1802 1305 1814
rect 1247 1742 1259 1802
rect 1293 1742 1305 1802
rect 1247 1730 1305 1742
rect 1376 1802 1434 1814
rect 1376 1742 1388 1802
rect 1422 1742 1434 1802
rect 1376 1730 1434 1742
rect 1465 1802 1522 1814
rect 1465 1742 1476 1802
rect 1510 1742 1522 1802
rect 1465 1730 1522 1742
rect 1552 1802 1610 1814
rect 1552 1742 1564 1802
rect 1598 1742 1610 1802
rect 1552 1730 1610 1742
rect 1682 1802 1740 1814
rect 1682 1742 1694 1802
rect 1728 1742 1740 1802
rect 1682 1730 1740 1742
rect 1770 1802 1828 1814
rect 1770 1742 1782 1802
rect 1816 1742 1828 1802
rect 1770 1730 1828 1742
rect 1858 1802 1916 1814
rect 1858 1742 1870 1802
rect 1904 1742 1916 1802
rect 1858 1730 1916 1742
rect 1988 1802 2046 1814
rect 1988 1742 2000 1802
rect 2034 1742 2046 1802
rect 1988 1730 2046 1742
rect 2076 1802 2134 1814
rect 2076 1742 2088 1802
rect 2122 1742 2134 1802
rect 2076 1730 2134 1742
rect 2206 1789 2264 1814
rect 2206 1755 2218 1789
rect 2252 1755 2264 1789
rect 2206 1730 2264 1755
rect 2294 1789 2352 1814
rect 2294 1755 2306 1789
rect 2340 1755 2352 1789
rect 2294 1730 2352 1755
rect 2382 1789 2440 1814
rect 2382 1755 2394 1789
rect 2428 1755 2440 1789
rect 2382 1730 2440 1755
rect 2624 1789 2682 1814
rect 2624 1755 2636 1789
rect 2670 1755 2682 1789
rect 2624 1730 2682 1755
rect 2712 1789 2770 1814
rect 2712 1755 2724 1789
rect 2758 1755 2770 1789
rect 2712 1730 2770 1755
rect 2954 1790 3012 1815
rect 2954 1756 2966 1790
rect 3000 1756 3012 1790
rect 2954 1731 3012 1756
rect 3042 1790 3100 1815
rect 3042 1756 3054 1790
rect 3088 1756 3100 1790
rect 3042 1731 3100 1756
rect 459 1216 517 1228
rect 459 1156 471 1216
rect 505 1156 517 1216
rect 459 1144 517 1156
rect 547 1216 605 1228
rect 547 1156 559 1216
rect 593 1156 605 1216
rect 547 1144 605 1156
rect 635 1216 693 1228
rect 635 1156 647 1216
rect 681 1156 693 1216
rect 635 1144 693 1156
rect 765 1216 823 1228
rect 765 1156 777 1216
rect 811 1156 823 1216
rect 765 1144 823 1156
rect 853 1216 911 1228
rect 853 1156 865 1216
rect 899 1156 911 1216
rect 853 1144 911 1156
rect 941 1216 999 1228
rect 941 1156 953 1216
rect 987 1156 999 1216
rect 941 1144 999 1156
rect 1071 1216 1129 1228
rect 1071 1156 1083 1216
rect 1117 1156 1129 1216
rect 1071 1144 1129 1156
rect 1159 1216 1217 1228
rect 1159 1156 1171 1216
rect 1205 1156 1217 1216
rect 1159 1144 1217 1156
rect 1247 1216 1305 1228
rect 1247 1156 1259 1216
rect 1293 1156 1305 1216
rect 1247 1144 1305 1156
rect 1376 1216 1434 1228
rect 1376 1156 1388 1216
rect 1422 1156 1434 1216
rect 1376 1144 1434 1156
rect 1465 1216 1522 1228
rect 1465 1156 1476 1216
rect 1510 1156 1522 1216
rect 1465 1144 1522 1156
rect 1552 1216 1610 1228
rect 1552 1156 1564 1216
rect 1598 1156 1610 1216
rect 1552 1144 1610 1156
rect 1682 1216 1740 1228
rect 1682 1156 1694 1216
rect 1728 1156 1740 1216
rect 1682 1144 1740 1156
rect 1770 1216 1828 1228
rect 1770 1156 1782 1216
rect 1816 1156 1828 1216
rect 1770 1144 1828 1156
rect 1858 1216 1916 1228
rect 1858 1156 1870 1216
rect 1904 1156 1916 1216
rect 1858 1144 1916 1156
rect 1988 1216 2046 1228
rect 1988 1156 2000 1216
rect 2034 1156 2046 1216
rect 1988 1144 2046 1156
rect 2076 1216 2134 1228
rect 2076 1156 2088 1216
rect 2122 1156 2134 1216
rect 2076 1144 2134 1156
rect 2206 1203 2264 1228
rect 2206 1169 2218 1203
rect 2252 1169 2264 1203
rect 2206 1144 2264 1169
rect 2294 1203 2352 1228
rect 2294 1169 2306 1203
rect 2340 1169 2352 1203
rect 2294 1144 2352 1169
rect 2382 1203 2440 1228
rect 2382 1169 2394 1203
rect 2428 1169 2440 1203
rect 2382 1144 2440 1169
rect 2624 1203 2682 1228
rect 2624 1169 2636 1203
rect 2670 1169 2682 1203
rect 2624 1144 2682 1169
rect 2712 1203 2770 1228
rect 2712 1169 2724 1203
rect 2758 1169 2770 1203
rect 2712 1144 2770 1169
rect 2842 1216 2900 1228
rect 2842 1080 2854 1216
rect 2888 1080 2900 1216
rect 2842 1068 2900 1080
rect 2930 1216 2988 1228
rect 2930 1080 2942 1216
rect 2976 1080 2988 1216
rect 2930 1068 2988 1080
rect 3060 1216 3118 1228
rect 3060 1080 3072 1216
rect 3106 1080 3118 1216
rect 3060 1068 3118 1080
rect 3148 1216 3206 1228
rect 3148 1080 3160 1216
rect 3194 1080 3206 1216
rect 3148 1068 3206 1080
rect 3278 1140 3336 1152
rect 3278 1080 3290 1140
rect 3324 1080 3336 1140
rect 3278 1068 3336 1080
rect 3366 1140 3424 1152
rect 3366 1080 3378 1140
rect 3412 1080 3424 1140
rect 3366 1068 3424 1080
rect 476 471 534 496
rect 476 437 488 471
rect 522 437 534 471
rect 476 412 534 437
rect 564 471 622 496
rect 564 437 576 471
rect 610 437 622 471
rect 564 412 622 437
rect 834 471 892 496
rect 834 437 846 471
rect 880 437 892 471
rect 834 412 892 437
rect 922 471 980 496
rect 922 437 934 471
rect 968 437 980 471
rect 922 412 980 437
rect 1010 471 1068 496
rect 1010 437 1022 471
rect 1056 437 1068 471
rect 1010 412 1068 437
rect 1412 484 1470 496
rect 1412 424 1424 484
rect 1458 424 1470 484
rect 1412 412 1470 424
rect 1500 484 1558 496
rect 1500 424 1512 484
rect 1546 424 1558 484
rect 1500 412 1558 424
rect 1588 484 1646 496
rect 1588 424 1600 484
rect 1634 424 1646 484
rect 1588 412 1646 424
rect 1883 471 1941 496
rect 1883 437 1895 471
rect 1929 437 1941 471
rect 1883 412 1941 437
rect 1971 471 2029 496
rect 1971 437 1983 471
rect 2017 437 2029 471
rect 1971 412 2029 437
rect 2244 471 2302 496
rect 2244 437 2256 471
rect 2290 437 2302 471
rect 2244 412 2302 437
rect 2332 471 2390 496
rect 2332 437 2344 471
rect 2378 437 2390 471
rect 2332 412 2390 437
rect 2420 471 2478 496
rect 2420 437 2432 471
rect 2466 437 2478 471
rect 2420 412 2478 437
rect 2508 471 2566 496
rect 2508 437 2520 471
rect 2554 437 2566 471
rect 2508 412 2566 437
rect 1456 271 1514 283
rect 1456 211 1468 271
rect 1502 211 1514 271
rect 1456 199 1514 211
rect 1544 271 1602 283
rect 1544 211 1556 271
rect 1590 211 1602 271
rect 1544 199 1602 211
rect 2750 471 2808 496
rect 2750 437 2762 471
rect 2796 437 2808 471
rect 2750 412 2808 437
rect 2838 471 2896 496
rect 2838 437 2850 471
rect 2884 437 2896 471
rect 2838 412 2896 437
rect 3119 471 3177 496
rect 3119 437 3131 471
rect 3165 437 3177 471
rect 3119 412 3177 437
rect 3207 471 3265 496
rect 3207 437 3219 471
rect 3253 437 3265 471
rect 3207 412 3265 437
rect 3295 471 3353 496
rect 3295 437 3307 471
rect 3341 437 3353 471
rect 3295 412 3353 437
rect 3537 471 3595 496
rect 3537 437 3549 471
rect 3583 437 3595 471
rect 3537 412 3595 437
rect 3625 471 3683 496
rect 3625 437 3637 471
rect 3671 437 3683 471
rect 3625 412 3683 437
<< ndiffc >>
rect 160 1406 194 1440
rect 248 1406 282 1440
rect 471 1393 505 1453
rect 559 1393 593 1453
rect 647 1393 681 1453
rect 777 1393 811 1453
rect 865 1393 899 1453
rect 953 1393 987 1453
rect 1083 1393 1117 1453
rect 1171 1393 1205 1453
rect 1259 1393 1293 1453
rect 1388 1393 1422 1453
rect 1476 1393 1510 1453
rect 1564 1393 1598 1453
rect 1694 1393 1728 1453
rect 1782 1393 1816 1453
rect 1870 1393 1904 1453
rect 2000 1393 2034 1453
rect 2088 1393 2122 1453
rect 2218 1406 2252 1440
rect 2306 1406 2340 1440
rect 2394 1406 2428 1440
rect 2636 1406 2670 1440
rect 2724 1406 2758 1440
rect 2966 1407 3000 1441
rect 3054 1407 3088 1441
rect 471 807 505 867
rect 559 807 593 867
rect 647 807 681 867
rect 777 807 811 867
rect 865 807 899 867
rect 953 807 987 867
rect 1083 807 1117 867
rect 1171 807 1205 867
rect 1259 807 1293 867
rect 1388 807 1422 867
rect 1476 807 1510 867
rect 1564 807 1598 867
rect 1694 807 1728 867
rect 1782 807 1816 867
rect 1870 807 1904 867
rect 2000 807 2034 867
rect 2088 807 2122 867
rect 2218 820 2252 854
rect 2306 820 2340 854
rect 2394 820 2428 854
rect 2636 820 2670 854
rect 2724 820 2758 854
rect 2854 706 2888 842
rect 2942 706 2976 842
rect 3072 706 3106 842
rect 3160 706 3194 842
rect 3290 782 3324 842
rect 3378 782 3412 842
rect 3501 706 3535 842
rect 3589 706 3623 842
rect 488 88 522 122
rect 576 88 610 122
rect 846 88 880 122
rect 934 88 968 122
rect 1022 88 1056 122
rect 1895 88 1929 122
rect 1983 88 2017 122
rect 2256 88 2290 122
rect 2344 88 2378 122
rect 2432 88 2466 122
rect 2520 88 2554 122
rect 2762 88 2796 122
rect 2850 88 2884 122
rect 3131 88 3165 122
rect 3219 88 3253 122
rect 3307 88 3341 122
rect 3549 88 3583 122
rect 3637 88 3671 122
<< pdiffc >>
rect 160 1755 194 1789
rect 248 1755 282 1789
rect 471 1742 505 1802
rect 559 1742 593 1802
rect 647 1742 681 1802
rect 777 1742 811 1802
rect 865 1742 899 1802
rect 953 1742 987 1802
rect 1083 1742 1117 1802
rect 1171 1742 1205 1802
rect 1259 1742 1293 1802
rect 1388 1742 1422 1802
rect 1476 1742 1510 1802
rect 1564 1742 1598 1802
rect 1694 1742 1728 1802
rect 1782 1742 1816 1802
rect 1870 1742 1904 1802
rect 2000 1742 2034 1802
rect 2088 1742 2122 1802
rect 2218 1755 2252 1789
rect 2306 1755 2340 1789
rect 2394 1755 2428 1789
rect 2636 1755 2670 1789
rect 2724 1755 2758 1789
rect 2966 1756 3000 1790
rect 3054 1756 3088 1790
rect 471 1156 505 1216
rect 559 1156 593 1216
rect 647 1156 681 1216
rect 777 1156 811 1216
rect 865 1156 899 1216
rect 953 1156 987 1216
rect 1083 1156 1117 1216
rect 1171 1156 1205 1216
rect 1259 1156 1293 1216
rect 1388 1156 1422 1216
rect 1476 1156 1510 1216
rect 1564 1156 1598 1216
rect 1694 1156 1728 1216
rect 1782 1156 1816 1216
rect 1870 1156 1904 1216
rect 2000 1156 2034 1216
rect 2088 1156 2122 1216
rect 2218 1169 2252 1203
rect 2306 1169 2340 1203
rect 2394 1169 2428 1203
rect 2636 1169 2670 1203
rect 2724 1169 2758 1203
rect 2854 1080 2888 1216
rect 2942 1080 2976 1216
rect 3072 1080 3106 1216
rect 3160 1080 3194 1216
rect 3290 1080 3324 1140
rect 3378 1080 3412 1140
rect 488 437 522 471
rect 576 437 610 471
rect 846 437 880 471
rect 934 437 968 471
rect 1022 437 1056 471
rect 1424 424 1458 484
rect 1512 424 1546 484
rect 1600 424 1634 484
rect 1895 437 1929 471
rect 1983 437 2017 471
rect 2256 437 2290 471
rect 2344 437 2378 471
rect 2432 437 2466 471
rect 2520 437 2554 471
rect 1468 211 1502 271
rect 1556 211 1590 271
rect 2762 437 2796 471
rect 2850 437 2884 471
rect 3131 437 3165 471
rect 3219 437 3253 471
rect 3307 437 3341 471
rect 3549 437 3583 471
rect 3637 437 3671 471
<< psubdiff >>
rect 36 1440 94 1477
rect 36 1406 48 1440
rect 82 1406 94 1440
rect 36 1369 94 1406
rect 2512 1440 2570 1477
rect 2512 1406 2524 1440
rect 2558 1406 2570 1440
rect 2512 1369 2570 1406
rect 2842 1441 2900 1478
rect 2842 1407 2854 1441
rect 2888 1407 2900 1441
rect 2842 1370 2900 1407
rect 2512 854 2570 891
rect 2512 820 2524 854
rect 2558 820 2570 854
rect 2512 783 2570 820
rect 364 122 422 159
rect 364 88 376 122
rect 410 88 422 122
rect 364 51 422 88
rect 1771 122 1829 159
rect 1771 88 1783 122
rect 1817 88 1829 122
rect 1771 51 1829 88
rect 2638 122 2696 159
rect 2638 88 2650 122
rect 2684 88 2696 122
rect 2638 51 2696 88
rect 3425 122 3483 159
rect 3425 88 3437 122
rect 3471 88 3483 122
rect 3425 51 3483 88
<< nsubdiff >>
rect 36 1789 94 1826
rect 36 1755 48 1789
rect 82 1755 94 1789
rect 36 1718 94 1755
rect 2512 1789 2570 1826
rect 2512 1755 2524 1789
rect 2558 1755 2570 1789
rect 2512 1718 2570 1755
rect 2842 1790 2900 1827
rect 2842 1756 2854 1790
rect 2888 1756 2900 1790
rect 2842 1719 2900 1756
rect 2512 1203 2570 1240
rect 2512 1169 2524 1203
rect 2558 1169 2570 1203
rect 2512 1132 2570 1169
rect 364 471 422 508
rect 364 437 376 471
rect 410 437 422 471
rect 364 400 422 437
rect 1771 471 1829 508
rect 1771 437 1783 471
rect 1817 437 1829 471
rect 1771 400 1829 437
rect 2638 471 2696 508
rect 2638 437 2650 471
rect 2684 437 2696 471
rect 2638 400 2696 437
rect 3425 471 3483 508
rect 3425 437 3437 471
rect 3471 437 3483 471
rect 3425 400 3483 437
<< psubdiffcont >>
rect 48 1406 82 1440
rect 2524 1406 2558 1440
rect 2854 1407 2888 1441
rect 2524 820 2558 854
rect 376 88 410 122
rect 1783 88 1817 122
rect 2650 88 2684 122
rect 3437 88 3471 122
<< nsubdiffcont >>
rect 48 1755 82 1789
rect 2524 1755 2558 1789
rect 2854 1756 2888 1790
rect 2524 1169 2558 1203
rect 376 437 410 471
rect 1783 437 1817 471
rect 2650 437 2684 471
rect 3437 437 3471 471
<< poly >>
rect 206 1814 236 1840
rect 517 1814 547 1840
rect 605 1814 635 1840
rect 823 1814 853 1840
rect 911 1814 941 1840
rect 1129 1814 1159 1840
rect 1217 1814 1247 1840
rect 1434 1814 1465 1840
rect 1522 1814 1552 1840
rect 1740 1814 1770 1840
rect 1828 1814 1858 1840
rect 2046 1814 2076 1840
rect 2264 1814 2294 1840
rect 2352 1814 2382 1840
rect 2682 1814 2712 1840
rect 206 1640 236 1730
rect 145 1624 236 1640
rect 145 1590 161 1624
rect 195 1590 236 1624
rect 145 1574 236 1590
rect 386 1624 452 1640
rect 517 1624 547 1730
rect 386 1590 402 1624
rect 436 1590 547 1624
rect 605 1618 635 1730
rect 386 1574 452 1590
rect 206 1465 236 1574
rect 517 1465 547 1590
rect 589 1602 655 1618
rect 589 1568 605 1602
rect 639 1568 655 1602
rect 589 1552 655 1568
rect 697 1602 751 1618
rect 823 1602 853 1730
rect 697 1568 707 1602
rect 741 1568 853 1602
rect 697 1552 751 1568
rect 605 1465 635 1552
rect 823 1465 853 1568
rect 911 1465 941 1730
rect 1003 1602 1057 1618
rect 1129 1602 1159 1730
rect 1003 1568 1013 1602
rect 1047 1568 1159 1602
rect 1003 1552 1057 1568
rect 1129 1465 1159 1568
rect 1217 1465 1247 1730
rect 1434 1704 1465 1730
rect 1309 1602 1363 1618
rect 1435 1602 1465 1704
rect 1309 1568 1319 1602
rect 1353 1568 1465 1602
rect 1309 1552 1363 1568
rect 1435 1491 1465 1568
rect 1434 1465 1465 1491
rect 1522 1465 1552 1730
rect 1614 1602 1668 1618
rect 1740 1602 1770 1730
rect 1614 1568 1624 1602
rect 1658 1568 1770 1602
rect 1614 1552 1668 1568
rect 1740 1465 1770 1568
rect 1828 1465 1858 1730
rect 1920 1602 1974 1618
rect 2046 1602 2076 1730
rect 2264 1698 2294 1730
rect 2214 1682 2294 1698
rect 2214 1648 2230 1682
rect 2264 1648 2294 1682
rect 2214 1632 2294 1648
rect 1920 1568 1930 1602
rect 1964 1568 2076 1602
rect 1920 1552 1974 1568
rect 2046 1465 2076 1568
rect 2264 1465 2294 1632
rect 2352 1553 2382 1730
rect 3012 1815 3042 1841
rect 2682 1640 2712 1730
rect 3012 1641 3042 1731
rect 2621 1624 2712 1640
rect 2621 1590 2637 1624
rect 2671 1590 2712 1624
rect 2621 1574 2712 1590
rect 2951 1625 3042 1641
rect 2951 1591 2967 1625
rect 3001 1591 3042 1625
rect 2951 1575 3042 1591
rect 2352 1537 2432 1553
rect 2352 1503 2382 1537
rect 2416 1503 2432 1537
rect 2352 1487 2432 1503
rect 2352 1465 2382 1487
rect 2682 1465 2712 1574
rect 206 1226 236 1381
rect 517 1355 547 1381
rect 605 1355 635 1381
rect 823 1355 853 1381
rect 911 1355 941 1381
rect 1129 1355 1159 1381
rect 1217 1355 1247 1381
rect 1434 1355 1465 1381
rect 1522 1355 1552 1381
rect 1740 1355 1770 1381
rect 1828 1355 1858 1381
rect 2046 1355 2076 1381
rect 2264 1355 2294 1381
rect 2352 1355 2382 1381
rect 3012 1466 3042 1575
rect 2682 1355 2712 1381
rect 3012 1356 3042 1382
rect 2884 1309 2950 1325
rect 2884 1275 2900 1309
rect 2934 1275 2950 1309
rect 2884 1259 2950 1275
rect 517 1228 547 1254
rect 605 1228 635 1254
rect 823 1228 853 1254
rect 911 1228 941 1254
rect 1129 1228 1159 1254
rect 1217 1228 1247 1254
rect 1434 1228 1465 1254
rect 1522 1228 1552 1254
rect 1740 1228 1770 1254
rect 1828 1228 1858 1254
rect 2046 1228 2076 1254
rect 2264 1228 2294 1254
rect 2352 1228 2382 1254
rect 188 1210 254 1226
rect 188 1176 204 1210
rect 238 1176 254 1210
rect 188 1160 254 1176
rect 2682 1228 2712 1254
rect 2900 1228 2930 1259
rect 3118 1228 3148 1254
rect 386 1038 452 1054
rect 517 1038 547 1144
rect 386 1004 402 1038
rect 436 1004 547 1038
rect 605 1032 635 1144
rect 386 988 452 1004
rect 517 879 547 1004
rect 589 1016 655 1032
rect 589 982 605 1016
rect 639 982 655 1016
rect 589 966 655 982
rect 697 1016 751 1032
rect 823 1016 853 1144
rect 697 982 707 1016
rect 741 982 853 1016
rect 697 966 751 982
rect 605 879 635 966
rect 823 879 853 982
rect 911 879 941 1144
rect 1003 1016 1057 1032
rect 1129 1016 1159 1144
rect 1003 982 1013 1016
rect 1047 982 1159 1016
rect 1003 966 1057 982
rect 1129 879 1159 982
rect 1217 879 1247 1144
rect 1434 1118 1465 1144
rect 1309 1016 1363 1032
rect 1435 1016 1465 1118
rect 1309 982 1319 1016
rect 1353 982 1465 1016
rect 1309 966 1363 982
rect 1435 905 1465 982
rect 1434 879 1465 905
rect 1522 879 1552 1144
rect 1614 1016 1668 1032
rect 1740 1016 1770 1144
rect 1614 982 1624 1016
rect 1658 982 1770 1016
rect 1614 966 1668 982
rect 1740 879 1770 982
rect 1828 879 1858 1144
rect 1920 1016 1974 1032
rect 2046 1016 2076 1144
rect 2264 1112 2294 1144
rect 2214 1096 2294 1112
rect 2214 1062 2230 1096
rect 2264 1062 2294 1096
rect 2214 1046 2294 1062
rect 1920 982 1930 1016
rect 1964 982 2076 1016
rect 1920 966 1974 982
rect 2046 879 2076 982
rect 2264 879 2294 1046
rect 2352 967 2382 1144
rect 2682 1054 2712 1144
rect 3336 1152 3366 1178
rect 2621 1038 2712 1054
rect 2900 1042 2930 1068
rect 2621 1004 2637 1038
rect 2671 1004 2712 1038
rect 2621 988 2712 1004
rect 2352 951 2432 967
rect 2352 917 2382 951
rect 2416 917 2432 951
rect 2352 901 2432 917
rect 2352 879 2382 901
rect 2682 879 2712 988
rect 3118 976 3148 1068
rect 3336 976 3366 1068
rect 2850 960 2930 976
rect 2850 926 2866 960
rect 2900 926 2930 960
rect 2850 910 2930 926
rect 3057 960 3148 976
rect 3057 926 3073 960
rect 3107 926 3148 960
rect 3057 910 3148 926
rect 3275 960 3366 976
rect 3275 926 3291 960
rect 3325 926 3366 960
rect 3520 994 3586 1010
rect 3520 960 3536 994
rect 3570 960 3586 994
rect 3520 944 3586 960
rect 3275 910 3366 926
rect 517 769 547 795
rect 605 769 635 795
rect 823 769 853 795
rect 911 769 941 795
rect 1129 769 1159 795
rect 1217 769 1247 795
rect 1434 769 1465 795
rect 1522 769 1552 795
rect 1740 769 1770 795
rect 1828 769 1858 795
rect 2046 769 2076 795
rect 2264 769 2294 795
rect 2352 769 2382 795
rect 2900 854 2930 910
rect 3118 854 3148 910
rect 3336 854 3366 910
rect 3547 854 3577 944
rect 2682 769 2712 795
rect 3336 744 3366 770
rect 2900 668 2930 694
rect 3118 668 3148 694
rect 3547 668 3577 694
rect 534 496 564 522
rect 892 496 922 522
rect 980 496 1010 522
rect 1470 496 1500 522
rect 1558 496 1588 522
rect 1941 496 1971 522
rect 2302 496 2332 522
rect 2390 496 2420 522
rect 2478 496 2508 522
rect 534 322 564 412
rect 892 380 922 412
rect 473 306 564 322
rect 842 364 922 380
rect 842 330 858 364
rect 892 330 922 364
rect 842 314 922 330
rect 473 272 489 306
rect 523 272 564 306
rect 473 256 564 272
rect 534 147 564 256
rect 892 147 922 314
rect 980 235 1010 412
rect 1470 385 1500 412
rect 1558 385 1588 412
rect 2808 496 2838 522
rect 3177 496 3207 522
rect 3265 496 3295 522
rect 1470 365 1588 385
rect 1470 355 1512 365
rect 1496 331 1512 355
rect 1546 355 1588 365
rect 1546 331 1562 355
rect 1496 313 1562 331
rect 1941 322 1971 412
rect 2302 381 2332 412
rect 1514 283 1544 313
rect 1880 306 1971 322
rect 2252 365 2332 381
rect 2252 331 2268 365
rect 2302 331 2332 365
rect 2252 315 2332 331
rect 980 219 1060 235
rect 980 185 1010 219
rect 1044 185 1060 219
rect 1880 272 1896 306
rect 1930 272 1971 306
rect 1880 256 1971 272
rect 980 169 1060 185
rect 1514 173 1544 199
rect 980 147 1010 169
rect 1941 147 1971 256
rect 2302 147 2332 315
rect 2390 310 2420 412
rect 2378 294 2432 310
rect 2378 260 2388 294
rect 2422 260 2432 294
rect 2378 244 2432 260
rect 2390 147 2420 244
rect 2478 235 2508 412
rect 3595 496 3625 522
rect 2808 322 2838 412
rect 3177 380 3207 412
rect 2747 306 2838 322
rect 3127 364 3207 380
rect 3127 330 3143 364
rect 3177 330 3207 364
rect 3127 314 3207 330
rect 2747 272 2763 306
rect 2797 272 2838 306
rect 2747 256 2838 272
rect 2478 219 2558 235
rect 2478 185 2508 219
rect 2542 185 2558 219
rect 2478 169 2558 185
rect 2478 147 2508 169
rect 534 37 564 63
rect 892 37 922 63
rect 980 37 1010 63
rect 2808 147 2838 256
rect 3177 147 3207 314
rect 3265 235 3295 412
rect 3595 322 3625 412
rect 3534 306 3625 322
rect 3534 272 3550 306
rect 3584 272 3625 306
rect 3534 256 3625 272
rect 3265 219 3345 235
rect 3265 185 3295 219
rect 3329 185 3345 219
rect 3265 169 3345 185
rect 3265 147 3295 169
rect 1941 37 1971 63
rect 2302 37 2332 63
rect 2390 37 2420 63
rect 2478 37 2508 63
rect 3595 147 3625 256
rect 2808 37 2838 63
rect 3177 37 3207 63
rect 3265 37 3295 63
rect 3595 37 3625 63
<< polycont >>
rect 161 1590 195 1624
rect 402 1590 436 1624
rect 605 1568 639 1602
rect 707 1568 741 1602
rect 1013 1568 1047 1602
rect 1319 1568 1353 1602
rect 1624 1568 1658 1602
rect 2230 1648 2264 1682
rect 1930 1568 1964 1602
rect 2637 1590 2671 1624
rect 2967 1591 3001 1625
rect 2382 1503 2416 1537
rect 2900 1275 2934 1309
rect 204 1176 238 1210
rect 402 1004 436 1038
rect 605 982 639 1016
rect 707 982 741 1016
rect 1013 982 1047 1016
rect 1319 982 1353 1016
rect 1624 982 1658 1016
rect 2230 1062 2264 1096
rect 1930 982 1964 1016
rect 2637 1004 2671 1038
rect 2382 917 2416 951
rect 2866 926 2900 960
rect 3073 926 3107 960
rect 3291 926 3325 960
rect 3536 960 3570 994
rect 858 330 892 364
rect 489 272 523 306
rect 1512 331 1546 365
rect 2268 331 2302 365
rect 1010 185 1044 219
rect 1896 272 1930 306
rect 2388 260 2422 294
rect 3143 330 3177 364
rect 2763 272 2797 306
rect 2508 185 2542 219
rect 3550 272 3584 306
rect 3295 185 3329 219
<< locali >>
rect 36 1789 194 1818
rect 36 1755 48 1789
rect 82 1755 160 1789
rect 36 1726 194 1755
rect 248 1789 282 1818
rect 248 1624 282 1755
rect 471 1802 505 1818
rect 145 1590 161 1624
rect 195 1590 211 1624
rect 48 1440 194 1469
rect 82 1406 160 1440
rect 48 1377 194 1406
rect 248 1440 282 1590
rect 402 1624 436 1640
rect 402 1574 436 1590
rect 471 1602 505 1742
rect 559 1802 593 1818
rect 559 1726 593 1742
rect 647 1802 681 1818
rect 777 1802 811 1818
rect 681 1742 741 1760
rect 647 1726 741 1742
rect 707 1602 741 1726
rect 248 1377 282 1406
rect 471 1568 605 1602
rect 639 1568 655 1602
rect 471 1453 505 1568
rect 707 1469 741 1568
rect 471 1377 505 1393
rect 559 1453 593 1469
rect 559 1377 593 1393
rect 647 1453 741 1469
rect 681 1435 741 1453
rect 777 1453 811 1742
rect 865 1802 899 1818
rect 865 1726 899 1742
rect 953 1802 987 1818
rect 1083 1802 1117 1818
rect 987 1742 1047 1760
rect 953 1726 1047 1742
rect 1013 1602 1047 1726
rect 1013 1469 1047 1568
rect 647 1377 681 1393
rect 777 1377 811 1393
rect 865 1453 899 1469
rect 865 1377 899 1393
rect 953 1453 1047 1469
rect 987 1435 1047 1453
rect 1083 1453 1117 1742
rect 1171 1802 1205 1818
rect 1171 1726 1205 1742
rect 1259 1802 1293 1818
rect 1388 1802 1422 1818
rect 1293 1742 1353 1760
rect 1259 1726 1353 1742
rect 1319 1602 1353 1726
rect 1319 1469 1353 1568
rect 953 1377 987 1393
rect 1083 1377 1117 1393
rect 1171 1453 1205 1469
rect 1171 1377 1205 1393
rect 1259 1453 1353 1469
rect 1293 1435 1353 1453
rect 1388 1453 1422 1742
rect 1476 1802 1510 1818
rect 1476 1726 1510 1742
rect 1564 1802 1598 1818
rect 1694 1802 1728 1818
rect 1598 1742 1658 1760
rect 1564 1726 1658 1742
rect 1624 1602 1658 1726
rect 1624 1469 1658 1568
rect 1259 1377 1293 1393
rect 1388 1377 1422 1393
rect 1476 1453 1510 1469
rect 1476 1377 1510 1393
rect 1564 1453 1658 1469
rect 1598 1435 1658 1453
rect 1694 1453 1728 1742
rect 1782 1802 1816 1818
rect 1782 1726 1816 1742
rect 1870 1802 1904 1818
rect 2000 1802 2034 1818
rect 1904 1742 1964 1760
rect 1870 1726 1964 1742
rect 2000 1726 2034 1742
rect 2088 1802 2122 1818
rect 1930 1602 1964 1726
rect 1930 1469 1964 1568
rect 2088 1537 2122 1742
rect 2218 1789 2252 1818
rect 2218 1726 2252 1755
rect 2306 1789 2340 1818
rect 2306 1726 2340 1755
rect 2394 1789 2428 1818
rect 2394 1726 2428 1755
rect 2512 1789 2670 1818
rect 2512 1755 2524 1789
rect 2558 1755 2636 1789
rect 2512 1726 2670 1755
rect 2724 1789 2758 1818
rect 2214 1648 2230 1682
rect 2264 1648 2280 1682
rect 2724 1624 2758 1755
rect 2842 1790 3000 1819
rect 2842 1756 2854 1790
rect 2888 1756 2966 1790
rect 2842 1727 3000 1756
rect 3054 1790 3088 1819
rect 3054 1625 3088 1756
rect 2621 1590 2637 1624
rect 2671 1590 2687 1624
rect 2951 1591 2967 1625
rect 3001 1591 3017 1625
rect 2218 1503 2230 1537
rect 2264 1503 2382 1537
rect 2416 1503 2432 1537
rect 1564 1377 1598 1393
rect 1694 1377 1728 1393
rect 1782 1453 1816 1469
rect 1782 1377 1816 1393
rect 1870 1453 1964 1469
rect 1904 1435 1964 1453
rect 2000 1453 2034 1469
rect 1870 1377 1904 1393
rect 2000 1377 2034 1393
rect 2088 1453 2122 1503
rect 2088 1377 2122 1393
rect 2218 1440 2252 1469
rect 2218 1377 2252 1406
rect 2306 1440 2340 1469
rect 2306 1377 2340 1406
rect 2394 1440 2428 1469
rect 2394 1377 2428 1406
rect 2524 1440 2670 1469
rect 2558 1406 2636 1440
rect 2524 1377 2670 1406
rect 2724 1440 2758 1590
rect 2724 1377 2758 1406
rect 2854 1441 3000 1470
rect 2888 1407 2966 1441
rect 2854 1378 3000 1407
rect 3054 1441 3088 1591
rect 3054 1309 3088 1407
rect 2884 1275 2900 1309
rect 2934 1275 3570 1309
rect 471 1216 505 1232
rect 188 1176 204 1210
rect 238 1176 436 1210
rect 402 1038 436 1176
rect 402 988 436 1004
rect 471 1016 505 1156
rect 559 1216 593 1232
rect 559 1140 593 1156
rect 647 1216 681 1232
rect 777 1216 811 1232
rect 681 1156 741 1174
rect 647 1140 741 1156
rect 707 1016 741 1140
rect 471 982 605 1016
rect 639 982 655 1016
rect 471 867 505 982
rect 707 883 741 982
rect 471 791 505 807
rect 559 867 593 883
rect 559 791 593 807
rect 647 867 741 883
rect 681 849 741 867
rect 777 867 811 1156
rect 865 1216 899 1232
rect 865 1140 899 1156
rect 953 1216 987 1232
rect 1083 1216 1117 1232
rect 987 1156 1047 1174
rect 953 1140 1047 1156
rect 1013 1016 1047 1140
rect 1013 883 1047 982
rect 647 791 681 807
rect 777 791 811 807
rect 865 867 899 883
rect 865 791 899 807
rect 953 867 1047 883
rect 987 849 1047 867
rect 1083 867 1117 1156
rect 1171 1216 1205 1232
rect 1171 1140 1205 1156
rect 1259 1216 1293 1232
rect 1388 1216 1422 1232
rect 1293 1156 1353 1174
rect 1259 1140 1353 1156
rect 1319 1016 1353 1140
rect 1319 883 1353 982
rect 953 791 987 807
rect 1083 791 1117 807
rect 1171 867 1205 883
rect 1171 791 1205 807
rect 1259 867 1353 883
rect 1293 849 1353 867
rect 1388 867 1422 1156
rect 1476 1216 1510 1232
rect 1476 1140 1510 1156
rect 1564 1216 1598 1232
rect 1694 1216 1728 1232
rect 1598 1156 1658 1174
rect 1564 1140 1658 1156
rect 1624 1016 1658 1140
rect 1624 883 1658 982
rect 1259 791 1293 807
rect 1388 791 1422 807
rect 1476 867 1510 883
rect 1476 791 1510 807
rect 1564 867 1658 883
rect 1598 849 1658 867
rect 1694 867 1728 1156
rect 1782 1216 1816 1232
rect 1782 1140 1816 1156
rect 1870 1216 1904 1232
rect 2000 1216 2034 1232
rect 1904 1156 1964 1174
rect 1870 1140 1964 1156
rect 2000 1140 2034 1156
rect 2088 1216 2122 1232
rect 1930 1016 1964 1140
rect 1930 883 1964 982
rect 2088 951 2122 1156
rect 2218 1203 2252 1232
rect 2218 1140 2252 1169
rect 2306 1203 2340 1232
rect 2306 1140 2340 1169
rect 2394 1203 2428 1232
rect 2394 1140 2428 1169
rect 2512 1203 2670 1232
rect 2512 1169 2524 1203
rect 2558 1169 2636 1203
rect 2512 1140 2670 1169
rect 2724 1203 2758 1232
rect 2214 1062 2230 1096
rect 2264 1062 2280 1096
rect 2724 1038 2758 1169
rect 2854 1216 2888 1232
rect 2854 1064 2888 1080
rect 2942 1216 2976 1232
rect 2621 1004 2637 1038
rect 2671 1004 2687 1038
rect 2218 917 2230 951
rect 2264 917 2382 951
rect 2416 917 2432 951
rect 1564 791 1598 807
rect 1694 791 1728 807
rect 1782 867 1816 883
rect 1782 791 1816 807
rect 1870 867 1964 883
rect 1904 849 1964 867
rect 2000 867 2034 883
rect 1870 791 1904 807
rect 2000 791 2034 807
rect 2088 867 2122 917
rect 2088 791 2122 807
rect 2218 854 2252 883
rect 2218 791 2252 820
rect 2306 854 2340 883
rect 2306 791 2340 820
rect 2394 854 2428 883
rect 2394 791 2428 820
rect 2524 854 2670 883
rect 2558 820 2636 854
rect 2524 791 2670 820
rect 2724 854 2758 1004
rect 2866 960 2900 976
rect 2866 910 2900 926
rect 2942 960 2976 1080
rect 3072 1216 3106 1232
rect 3072 1064 3106 1080
rect 3160 1216 3194 1232
rect 3160 960 3194 1080
rect 3290 1140 3324 1156
rect 3290 1064 3324 1080
rect 3378 1140 3412 1156
rect 2942 926 3073 960
rect 3107 926 3123 960
rect 3160 926 3291 960
rect 3325 926 3341 960
rect 2724 791 2758 820
rect 2854 842 2888 858
rect 2854 690 2888 706
rect 2942 842 2976 926
rect 2942 690 2976 706
rect 3072 842 3106 858
rect 3072 690 3106 706
rect 3160 842 3194 926
rect 3378 888 3412 1080
rect 3536 994 3570 1275
rect 3536 944 3570 960
rect 3290 842 3324 858
rect 3290 766 3324 782
rect 3378 854 3535 888
rect 3378 842 3412 854
rect 3378 766 3412 782
rect 3501 842 3535 854
rect 364 471 522 500
rect 364 437 376 471
rect 410 437 488 471
rect 364 408 522 437
rect 576 471 610 500
rect 576 306 610 437
rect 846 471 880 500
rect 846 408 880 437
rect 934 471 968 500
rect 934 408 968 437
rect 1022 471 1056 500
rect 1022 408 1056 437
rect 1424 484 1458 614
rect 842 330 858 364
rect 892 330 908 364
rect 473 272 489 306
rect 523 272 539 306
rect 376 122 522 151
rect 410 88 488 122
rect 376 59 522 88
rect 576 122 610 272
rect 1424 292 1458 424
rect 1512 484 1546 500
rect 1512 408 1546 424
rect 1600 484 1634 615
rect 3160 602 3194 706
rect 3501 690 3535 706
rect 3589 842 3623 858
rect 3589 690 3623 706
rect 3049 568 3194 602
rect 1496 331 1512 365
rect 1546 331 1562 365
rect 1600 292 1634 424
rect 1771 471 1929 500
rect 1771 437 1783 471
rect 1817 437 1895 471
rect 1771 408 1929 437
rect 1983 471 2017 500
rect 1983 306 2017 437
rect 2256 471 2290 500
rect 2256 408 2290 437
rect 2344 471 2378 500
rect 2344 408 2378 437
rect 2432 471 2466 500
rect 2432 408 2466 437
rect 2520 471 2554 500
rect 2520 408 2554 437
rect 2638 471 2796 500
rect 2638 437 2650 471
rect 2684 437 2762 471
rect 2638 408 2796 437
rect 2850 471 2884 500
rect 2252 331 2268 365
rect 2302 331 2318 365
rect 2850 306 2884 437
rect 3049 364 3083 568
rect 3131 471 3165 500
rect 3131 408 3165 437
rect 3219 471 3253 500
rect 3219 408 3253 437
rect 3307 471 3341 500
rect 3307 408 3341 437
rect 3425 471 3583 500
rect 3425 437 3437 471
rect 3471 437 3549 471
rect 3425 408 3583 437
rect 3637 471 3671 500
rect 3049 330 3143 364
rect 3177 330 3193 364
rect 3637 306 3671 437
rect 1424 291 1468 292
rect 1590 291 1634 292
rect 1424 271 1502 291
rect 1424 257 1468 271
rect 846 185 858 219
rect 892 185 1010 219
rect 1044 185 1060 219
rect 1468 195 1502 211
rect 1556 271 1634 291
rect 1880 272 1896 306
rect 1930 272 1946 306
rect 1590 257 1634 271
rect 1556 195 1590 211
rect 576 59 610 88
rect 846 122 880 151
rect 846 59 880 88
rect 934 122 968 151
rect 934 59 968 88
rect 1022 122 1056 151
rect 1022 59 1056 88
rect 1783 122 1929 151
rect 1817 88 1895 122
rect 1783 59 1929 88
rect 1983 122 2017 272
rect 2372 260 2388 294
rect 2422 260 2438 294
rect 2747 272 2763 306
rect 2797 272 2813 306
rect 3534 272 3550 306
rect 3584 272 3600 306
rect 2372 185 2388 219
rect 2422 185 2508 219
rect 2542 185 2645 219
rect 1983 59 2017 88
rect 2256 122 2290 151
rect 2256 59 2290 88
rect 2344 122 2378 151
rect 2344 59 2378 88
rect 2432 122 2466 151
rect 2432 59 2466 88
rect 2520 122 2554 151
rect 2520 59 2554 88
rect 2650 122 2796 151
rect 2684 88 2762 122
rect 2650 59 2796 88
rect 2850 122 2884 272
rect 3131 185 3143 219
rect 3177 185 3295 219
rect 3329 185 3345 219
rect 2850 59 2884 88
rect 3131 122 3165 151
rect 3131 59 3165 88
rect 3219 122 3253 151
rect 3219 59 3253 88
rect 3307 122 3341 151
rect 3307 59 3341 88
rect 3437 122 3583 151
rect 3471 88 3549 122
rect 3437 59 3583 88
rect 3637 122 3671 272
rect 3637 59 3671 88
<< viali >>
rect 160 1755 194 1789
rect 248 1755 282 1789
rect 471 1742 505 1802
rect 161 1590 195 1624
rect 248 1590 282 1624
rect 160 1406 194 1440
rect 402 1590 436 1624
rect 559 1742 593 1802
rect 647 1742 681 1802
rect 248 1406 282 1440
rect 471 1393 505 1453
rect 559 1393 593 1453
rect 647 1393 681 1453
rect 777 1742 811 1802
rect 865 1742 899 1802
rect 953 1742 987 1802
rect 777 1393 811 1453
rect 865 1393 899 1453
rect 953 1393 987 1453
rect 1083 1742 1117 1802
rect 1171 1742 1205 1802
rect 1259 1742 1293 1802
rect 1083 1393 1117 1453
rect 1171 1393 1205 1453
rect 1259 1393 1293 1453
rect 1388 1742 1422 1802
rect 1476 1742 1510 1802
rect 1564 1742 1598 1802
rect 1388 1393 1422 1453
rect 1476 1393 1510 1453
rect 1564 1393 1598 1453
rect 1694 1742 1728 1802
rect 1782 1742 1816 1802
rect 1870 1742 1904 1802
rect 2000 1742 2034 1802
rect 2088 1742 2122 1802
rect 2218 1755 2252 1789
rect 2306 1755 2340 1789
rect 2394 1755 2428 1789
rect 2636 1755 2670 1789
rect 2724 1755 2758 1789
rect 2230 1648 2264 1682
rect 2966 1756 3000 1790
rect 3054 1756 3088 1790
rect 2637 1590 2671 1624
rect 2724 1590 2758 1624
rect 2967 1591 3001 1625
rect 3054 1591 3088 1625
rect 2088 1503 2122 1537
rect 2230 1503 2264 1537
rect 1694 1393 1728 1453
rect 1782 1393 1816 1453
rect 1870 1393 1904 1453
rect 2000 1393 2034 1453
rect 2088 1393 2122 1453
rect 2218 1406 2252 1440
rect 2306 1406 2340 1440
rect 2394 1406 2428 1440
rect 2636 1406 2670 1440
rect 2724 1406 2758 1440
rect 2966 1407 3000 1441
rect 3054 1407 3088 1441
rect 402 1004 436 1038
rect 471 1156 505 1216
rect 559 1156 593 1216
rect 647 1156 681 1216
rect 471 807 505 867
rect 559 807 593 867
rect 647 807 681 867
rect 777 1156 811 1216
rect 865 1156 899 1216
rect 953 1156 987 1216
rect 777 807 811 867
rect 865 807 899 867
rect 953 807 987 867
rect 1083 1156 1117 1216
rect 1171 1156 1205 1216
rect 1259 1156 1293 1216
rect 1083 807 1117 867
rect 1171 807 1205 867
rect 1259 807 1293 867
rect 1388 1156 1422 1216
rect 1476 1156 1510 1216
rect 1564 1156 1598 1216
rect 1388 807 1422 867
rect 1476 807 1510 867
rect 1564 807 1598 867
rect 1694 1156 1728 1216
rect 1782 1156 1816 1216
rect 1870 1156 1904 1216
rect 2000 1156 2034 1216
rect 2088 1156 2122 1216
rect 2218 1169 2252 1203
rect 2306 1169 2340 1203
rect 2394 1169 2428 1203
rect 2636 1169 2670 1203
rect 2724 1169 2758 1203
rect 2230 1062 2264 1096
rect 2854 1080 2888 1216
rect 2942 1080 2976 1216
rect 2637 1004 2671 1038
rect 2724 1004 2758 1038
rect 2088 917 2122 951
rect 2230 917 2264 951
rect 1694 807 1728 867
rect 1782 807 1816 867
rect 1870 807 1904 867
rect 2000 807 2034 867
rect 2088 807 2122 867
rect 2218 820 2252 854
rect 2306 820 2340 854
rect 2394 820 2428 854
rect 2636 820 2670 854
rect 2866 926 2900 960
rect 3072 1080 3106 1216
rect 3160 1080 3194 1216
rect 3290 1080 3324 1140
rect 3378 1080 3412 1140
rect 2724 820 2758 854
rect 2854 706 2888 842
rect 2942 706 2976 842
rect 3072 706 3106 842
rect 3160 706 3194 842
rect 3290 782 3324 842
rect 3378 782 3412 842
rect 1424 614 1458 648
rect 488 437 522 471
rect 576 437 610 471
rect 846 437 880 471
rect 934 437 968 471
rect 1022 437 1056 471
rect 1600 615 1634 649
rect 1424 424 1458 484
rect 858 330 892 364
rect 489 272 523 306
rect 576 272 610 306
rect 488 88 522 122
rect 1512 424 1546 484
rect 3501 706 3535 842
rect 3589 706 3623 842
rect 1600 424 1634 484
rect 1512 331 1546 365
rect 1895 437 1929 471
rect 1983 437 2017 471
rect 2256 437 2290 471
rect 2344 437 2378 471
rect 2432 437 2466 471
rect 2520 437 2554 471
rect 2762 437 2796 471
rect 2850 437 2884 471
rect 2268 331 2302 365
rect 3131 437 3165 471
rect 3219 437 3253 471
rect 3307 437 3341 471
rect 3549 437 3583 471
rect 3637 437 3671 471
rect 3143 330 3177 364
rect 858 185 892 219
rect 1468 211 1502 271
rect 1896 272 1930 306
rect 1983 272 2017 306
rect 1556 211 1590 271
rect 576 88 610 122
rect 846 88 880 122
rect 934 88 968 122
rect 1022 88 1056 122
rect 1895 88 1929 122
rect 2388 260 2422 294
rect 2763 272 2797 306
rect 2850 272 2884 306
rect 3550 272 3584 306
rect 3637 272 3671 306
rect 2388 185 2422 219
rect 2645 185 2679 219
rect 1983 88 2017 122
rect 2256 88 2290 122
rect 2344 88 2378 122
rect 2432 88 2466 122
rect 2520 88 2554 122
rect 2762 88 2796 122
rect 3143 185 3177 219
rect 2850 88 2884 122
rect 3131 88 3165 122
rect 3219 88 3253 122
rect 3307 88 3341 122
rect 3549 88 3583 122
rect 3637 88 3671 122
<< metal1 >>
rect 2467 2425 2477 2477
rect 2529 2425 2539 2477
rect 2487 2011 2521 2425
rect 2467 1959 2477 2011
rect 2530 1959 2540 2011
rect 2806 1876 3136 1877
rect 0 1843 3136 1876
rect 0 1842 2806 1843
rect 160 1814 194 1842
rect 154 1789 200 1814
rect 154 1755 160 1789
rect 194 1755 200 1789
rect 154 1730 200 1755
rect 242 1789 288 1814
rect 340 1789 350 1842
rect 402 1789 412 1842
rect 559 1814 593 1842
rect 865 1814 899 1842
rect 1170 1814 1204 1842
rect 1476 1814 1510 1842
rect 1782 1814 1816 1842
rect 2000 1814 2034 1842
rect 2218 1814 2252 1842
rect 2394 1814 2428 1842
rect 2636 1814 2670 1842
rect 2966 1815 3000 1843
rect 465 1802 511 1814
rect 242 1755 248 1789
rect 282 1755 288 1789
rect 242 1730 288 1755
rect 465 1742 471 1802
rect 505 1742 511 1802
rect 465 1730 511 1742
rect 553 1802 599 1814
rect 553 1742 559 1802
rect 593 1742 599 1802
rect 553 1730 599 1742
rect 641 1802 687 1814
rect 641 1742 647 1802
rect 681 1742 687 1802
rect 641 1730 687 1742
rect 771 1802 817 1814
rect 771 1742 777 1802
rect 811 1742 817 1802
rect 771 1730 817 1742
rect 859 1802 905 1814
rect 859 1742 865 1802
rect 899 1742 905 1802
rect 859 1730 905 1742
rect 947 1802 993 1814
rect 947 1742 953 1802
rect 987 1742 993 1802
rect 947 1730 993 1742
rect 1077 1802 1123 1814
rect 1077 1742 1083 1802
rect 1117 1742 1123 1802
rect 1077 1730 1123 1742
rect 1165 1802 1211 1814
rect 1165 1742 1171 1802
rect 1205 1742 1211 1802
rect 1165 1730 1211 1742
rect 1253 1802 1299 1814
rect 1253 1742 1259 1802
rect 1293 1742 1299 1802
rect 1253 1730 1299 1742
rect 1382 1802 1428 1814
rect 1382 1742 1388 1802
rect 1422 1742 1428 1802
rect 1382 1730 1428 1742
rect 1470 1802 1516 1814
rect 1470 1742 1476 1802
rect 1510 1742 1516 1802
rect 1470 1730 1516 1742
rect 1558 1802 1604 1814
rect 1558 1742 1564 1802
rect 1598 1742 1604 1802
rect 1558 1730 1604 1742
rect 1688 1802 1734 1814
rect 1688 1742 1694 1802
rect 1728 1742 1734 1802
rect 1688 1730 1734 1742
rect 1776 1802 1822 1814
rect 1776 1742 1782 1802
rect 1816 1742 1822 1802
rect 1776 1730 1822 1742
rect 1864 1802 1910 1814
rect 1864 1742 1870 1802
rect 1904 1742 1910 1802
rect 1864 1730 1910 1742
rect 1994 1802 2040 1814
rect 1994 1742 2000 1802
rect 2034 1742 2040 1802
rect 1994 1730 2040 1742
rect 2082 1802 2128 1814
rect 2082 1742 2088 1802
rect 2122 1742 2128 1802
rect 2082 1730 2128 1742
rect 2212 1789 2258 1814
rect 2212 1755 2218 1789
rect 2252 1755 2258 1789
rect 2212 1730 2258 1755
rect 2300 1789 2346 1814
rect 2300 1755 2306 1789
rect 2340 1755 2346 1789
rect 2300 1730 2346 1755
rect 2388 1789 2434 1814
rect 2388 1755 2394 1789
rect 2428 1755 2434 1789
rect 2388 1730 2434 1755
rect 2630 1789 2676 1814
rect 2630 1755 2636 1789
rect 2670 1755 2676 1789
rect 2630 1730 2676 1755
rect 2718 1789 2764 1814
rect 2718 1755 2724 1789
rect 2758 1755 2764 1789
rect 2718 1730 2764 1755
rect 2960 1790 3006 1815
rect 2960 1756 2966 1790
rect 3000 1756 3006 1790
rect 2960 1731 3006 1756
rect 3048 1790 3094 1815
rect 3048 1756 3054 1790
rect 3088 1756 3094 1790
rect 3048 1731 3094 1756
rect 2218 1682 2276 1688
rect 635 1648 2230 1682
rect 2264 1648 2276 1682
rect 149 1624 207 1630
rect 0 1590 161 1624
rect 195 1590 207 1624
rect 149 1584 207 1590
rect 236 1624 294 1630
rect 390 1624 448 1630
rect 635 1624 663 1648
rect 2218 1642 2276 1648
rect 236 1590 248 1624
rect 282 1590 402 1624
rect 436 1590 663 1624
rect 2306 1624 2340 1730
rect 2625 1624 2683 1630
rect 2306 1590 2637 1624
rect 2671 1590 2683 1624
rect 236 1584 294 1590
rect 390 1584 448 1590
rect 2076 1537 2134 1543
rect 2218 1537 2276 1543
rect 2076 1503 2088 1537
rect 2122 1503 2230 1537
rect 2264 1503 2276 1537
rect 2076 1497 2134 1503
rect 2218 1497 2276 1503
rect 2394 1465 2428 1590
rect 2625 1584 2683 1590
rect 2712 1624 2770 1630
rect 2955 1625 3013 1631
rect 2806 1624 2967 1625
rect 2712 1590 2724 1624
rect 2758 1591 2967 1624
rect 3001 1591 3013 1625
rect 2758 1590 2806 1591
rect 2712 1584 2770 1590
rect 2955 1585 3013 1591
rect 3042 1625 3100 1631
rect 3042 1591 3054 1625
rect 3088 1591 3136 1625
rect 3042 1585 3100 1591
rect 154 1440 200 1465
rect 154 1406 160 1440
rect 194 1406 200 1440
rect 154 1381 200 1406
rect 242 1440 288 1465
rect 242 1406 248 1440
rect 282 1406 288 1440
rect 242 1381 288 1406
rect 465 1453 511 1465
rect 465 1393 471 1453
rect 505 1393 511 1453
rect 465 1381 511 1393
rect 553 1453 599 1465
rect 553 1393 559 1453
rect 593 1393 599 1453
rect 553 1381 599 1393
rect 641 1453 687 1465
rect 641 1393 647 1453
rect 681 1393 687 1453
rect 641 1381 687 1393
rect 771 1453 817 1465
rect 771 1393 777 1453
rect 811 1393 817 1453
rect 771 1381 817 1393
rect 859 1453 905 1465
rect 859 1393 865 1453
rect 899 1393 905 1453
rect 859 1381 905 1393
rect 947 1453 993 1465
rect 947 1393 953 1453
rect 987 1393 993 1453
rect 947 1381 993 1393
rect 1077 1453 1123 1465
rect 1077 1393 1083 1453
rect 1117 1393 1123 1453
rect 1077 1381 1123 1393
rect 1165 1453 1211 1465
rect 1165 1393 1171 1453
rect 1205 1393 1211 1453
rect 1165 1381 1211 1393
rect 1253 1453 1299 1465
rect 1253 1393 1259 1453
rect 1293 1393 1299 1453
rect 1253 1381 1299 1393
rect 1382 1453 1428 1465
rect 1382 1393 1388 1453
rect 1422 1393 1428 1453
rect 1382 1381 1428 1393
rect 1470 1453 1516 1465
rect 1470 1393 1476 1453
rect 1510 1393 1516 1453
rect 1470 1381 1516 1393
rect 1558 1453 1604 1465
rect 1558 1393 1564 1453
rect 1598 1393 1604 1453
rect 1558 1381 1604 1393
rect 1688 1453 1734 1465
rect 1688 1393 1694 1453
rect 1728 1393 1734 1453
rect 1688 1381 1734 1393
rect 1776 1453 1822 1465
rect 1776 1393 1782 1453
rect 1816 1393 1822 1453
rect 1776 1381 1822 1393
rect 1864 1453 1910 1465
rect 1864 1393 1870 1453
rect 1904 1393 1910 1453
rect 1864 1381 1910 1393
rect 1994 1453 2040 1465
rect 1994 1393 2000 1453
rect 2034 1393 2040 1453
rect 1994 1381 2040 1393
rect 2082 1453 2128 1465
rect 2082 1393 2088 1453
rect 2122 1393 2128 1453
rect 2082 1381 2128 1393
rect 2212 1440 2258 1465
rect 2212 1406 2218 1440
rect 2252 1406 2258 1440
rect 2212 1381 2258 1406
rect 2300 1440 2346 1465
rect 2300 1406 2306 1440
rect 2340 1406 2346 1440
rect 2300 1381 2346 1406
rect 2388 1440 2434 1465
rect 2388 1406 2394 1440
rect 2428 1406 2434 1440
rect 2388 1381 2434 1406
rect 2630 1440 2676 1465
rect 2630 1406 2636 1440
rect 2670 1406 2676 1440
rect 2630 1381 2676 1406
rect 2718 1440 2764 1465
rect 2718 1406 2724 1440
rect 2758 1406 2764 1440
rect 2718 1381 2764 1406
rect 2960 1441 3006 1466
rect 2960 1407 2966 1441
rect 3000 1407 3006 1441
rect 2960 1382 3006 1407
rect 3048 1441 3094 1466
rect 3048 1407 3054 1441
rect 3088 1407 3094 1441
rect 3048 1382 3094 1407
rect 160 1352 194 1381
rect 559 1352 593 1381
rect 865 1352 899 1381
rect 1171 1352 1205 1381
rect 1476 1352 1510 1381
rect 2000 1352 2034 1381
rect 2218 1352 2252 1381
rect 2636 1352 2670 1381
rect 2966 1353 3000 1382
rect 2806 1352 3704 1353
rect 0 1319 3704 1352
rect 0 1318 2806 1319
rect 2854 1290 3024 1291
rect 0 1256 3324 1290
rect 0 1255 350 1256
rect 340 1203 350 1255
rect 402 1203 412 1256
rect 559 1228 593 1256
rect 865 1228 899 1256
rect 1170 1228 1204 1256
rect 1476 1228 1510 1256
rect 1782 1228 1816 1256
rect 2000 1228 2034 1256
rect 2218 1228 2252 1256
rect 2394 1228 2428 1256
rect 2636 1228 2670 1256
rect 2854 1228 2888 1256
rect 3072 1228 3106 1256
rect 465 1216 511 1228
rect 465 1156 471 1216
rect 505 1156 511 1216
rect 465 1144 511 1156
rect 553 1216 599 1228
rect 553 1156 559 1216
rect 593 1156 599 1216
rect 553 1144 599 1156
rect 641 1216 687 1228
rect 641 1156 647 1216
rect 681 1156 687 1216
rect 641 1144 687 1156
rect 771 1216 817 1228
rect 771 1156 777 1216
rect 811 1156 817 1216
rect 771 1144 817 1156
rect 859 1216 905 1228
rect 859 1156 865 1216
rect 899 1156 905 1216
rect 859 1144 905 1156
rect 947 1216 993 1228
rect 947 1156 953 1216
rect 987 1156 993 1216
rect 947 1144 993 1156
rect 1077 1216 1123 1228
rect 1077 1156 1083 1216
rect 1117 1156 1123 1216
rect 1077 1144 1123 1156
rect 1165 1216 1211 1228
rect 1165 1156 1171 1216
rect 1205 1156 1211 1216
rect 1165 1144 1211 1156
rect 1253 1216 1299 1228
rect 1253 1156 1259 1216
rect 1293 1156 1299 1216
rect 1253 1144 1299 1156
rect 1382 1216 1428 1228
rect 1382 1156 1388 1216
rect 1422 1156 1428 1216
rect 1382 1144 1428 1156
rect 1470 1216 1516 1228
rect 1470 1156 1476 1216
rect 1510 1156 1516 1216
rect 1470 1144 1516 1156
rect 1558 1216 1604 1228
rect 1558 1156 1564 1216
rect 1598 1156 1604 1216
rect 1558 1144 1604 1156
rect 1688 1216 1734 1228
rect 1688 1156 1694 1216
rect 1728 1156 1734 1216
rect 1688 1144 1734 1156
rect 1776 1216 1822 1228
rect 1776 1156 1782 1216
rect 1816 1156 1822 1216
rect 1776 1144 1822 1156
rect 1864 1216 1910 1228
rect 1864 1156 1870 1216
rect 1904 1156 1910 1216
rect 1864 1144 1910 1156
rect 1994 1216 2040 1228
rect 1994 1156 2000 1216
rect 2034 1156 2040 1216
rect 1994 1144 2040 1156
rect 2082 1216 2128 1228
rect 2082 1156 2088 1216
rect 2122 1156 2128 1216
rect 2082 1144 2128 1156
rect 2212 1203 2258 1228
rect 2212 1169 2218 1203
rect 2252 1169 2258 1203
rect 2212 1144 2258 1169
rect 2300 1203 2346 1228
rect 2300 1169 2306 1203
rect 2340 1169 2346 1203
rect 2300 1144 2346 1169
rect 2388 1203 2434 1228
rect 2388 1169 2394 1203
rect 2428 1169 2434 1203
rect 2388 1144 2434 1169
rect 2630 1203 2676 1228
rect 2630 1169 2636 1203
rect 2670 1169 2676 1203
rect 2630 1144 2676 1169
rect 2718 1203 2764 1228
rect 2718 1169 2724 1203
rect 2758 1169 2764 1203
rect 2718 1144 2764 1169
rect 2848 1216 2894 1228
rect 2218 1096 2276 1102
rect 635 1062 2230 1096
rect 2264 1062 2276 1096
rect 390 1038 448 1044
rect 635 1038 663 1062
rect 2218 1056 2276 1062
rect 0 1035 145 1038
rect 0 1004 83 1035
rect 73 983 83 1004
rect 135 983 145 1035
rect 330 1004 402 1038
rect 436 1004 663 1038
rect 2306 1038 2340 1144
rect 2848 1080 2854 1216
rect 2888 1080 2894 1216
rect 2848 1068 2894 1080
rect 2936 1216 2982 1228
rect 2936 1080 2942 1216
rect 2976 1080 2982 1216
rect 2936 1068 2982 1080
rect 3066 1216 3112 1228
rect 3066 1080 3072 1216
rect 3106 1080 3112 1216
rect 3066 1068 3112 1080
rect 3154 1216 3200 1228
rect 3154 1080 3160 1216
rect 3194 1080 3200 1216
rect 3290 1152 3324 1256
rect 3154 1068 3200 1080
rect 3284 1140 3330 1152
rect 3284 1080 3290 1140
rect 3324 1080 3330 1140
rect 3284 1068 3330 1080
rect 3372 1140 3418 1152
rect 3372 1080 3378 1140
rect 3412 1080 3418 1140
rect 3372 1068 3418 1080
rect 2625 1038 2683 1044
rect 2306 1004 2637 1038
rect 2671 1004 2683 1038
rect 390 998 448 1004
rect 2076 951 2134 957
rect 2218 951 2276 957
rect 2076 917 2088 951
rect 2122 917 2230 951
rect 2264 917 2276 951
rect 2076 911 2134 917
rect 2218 911 2276 917
rect 2394 879 2428 1004
rect 2625 998 2683 1004
rect 2712 1038 2770 1044
rect 2712 1004 2724 1038
rect 2758 1004 2900 1038
rect 2712 998 2770 1004
rect 2866 966 2900 1004
rect 2854 960 2912 966
rect 2854 926 2866 960
rect 2900 926 3623 960
rect 2854 920 2912 926
rect 465 867 511 879
rect 465 807 471 867
rect 505 807 511 867
rect 465 795 511 807
rect 553 867 599 879
rect 553 807 559 867
rect 593 807 599 867
rect 553 795 599 807
rect 641 867 687 879
rect 641 807 647 867
rect 681 807 687 867
rect 641 795 687 807
rect 771 867 817 879
rect 771 807 777 867
rect 811 807 817 867
rect 771 795 817 807
rect 859 867 905 879
rect 859 807 865 867
rect 899 807 905 867
rect 859 795 905 807
rect 947 867 993 879
rect 947 807 953 867
rect 987 807 993 867
rect 947 795 993 807
rect 1077 867 1123 879
rect 1077 807 1083 867
rect 1117 807 1123 867
rect 1077 795 1123 807
rect 1165 867 1211 879
rect 1165 807 1171 867
rect 1205 807 1211 867
rect 1165 795 1211 807
rect 1253 867 1299 879
rect 1253 807 1259 867
rect 1293 807 1299 867
rect 1253 795 1299 807
rect 1382 867 1428 879
rect 1382 807 1388 867
rect 1422 807 1428 867
rect 1382 795 1428 807
rect 1470 867 1516 879
rect 1470 807 1476 867
rect 1510 807 1516 867
rect 1470 795 1516 807
rect 1558 867 1604 879
rect 1558 807 1564 867
rect 1598 807 1604 867
rect 1558 795 1604 807
rect 1688 867 1734 879
rect 1688 807 1694 867
rect 1728 807 1734 867
rect 1688 795 1734 807
rect 1776 867 1822 879
rect 1776 807 1782 867
rect 1816 807 1822 867
rect 1776 795 1822 807
rect 1864 867 1910 879
rect 1864 807 1870 867
rect 1904 807 1910 867
rect 1864 795 1910 807
rect 1994 867 2040 879
rect 1994 807 2000 867
rect 2034 807 2040 867
rect 1994 795 2040 807
rect 2082 867 2128 879
rect 2082 807 2088 867
rect 2122 807 2128 867
rect 2082 795 2128 807
rect 2212 854 2258 879
rect 2212 820 2218 854
rect 2252 820 2258 854
rect 2212 795 2258 820
rect 2300 854 2346 879
rect 2300 820 2306 854
rect 2340 820 2346 854
rect 2300 795 2346 820
rect 2388 854 2434 879
rect 2388 820 2394 854
rect 2428 820 2434 854
rect 2388 795 2434 820
rect 2630 854 2676 879
rect 2630 820 2636 854
rect 2670 820 2676 854
rect 2630 795 2676 820
rect 2718 854 2764 879
rect 3589 854 3623 926
rect 2718 820 2724 854
rect 2758 820 2764 854
rect 2718 795 2764 820
rect 2848 842 2894 854
rect 559 766 593 795
rect 865 766 899 795
rect 1171 766 1205 795
rect 1476 766 1510 795
rect 2000 766 2034 795
rect 2218 766 2252 795
rect 2636 766 2670 795
rect 2848 766 2854 842
rect 0 732 2854 766
rect 2848 706 2854 732
rect 2888 706 2894 842
rect 2848 694 2894 706
rect 2936 842 2982 854
rect 2936 706 2942 842
rect 2976 706 2982 842
rect 2936 694 2982 706
rect 3066 842 3112 854
rect 3066 706 3072 842
rect 3106 706 3112 842
rect 3066 694 3112 706
rect 3154 842 3200 854
rect 3154 706 3160 842
rect 3194 706 3200 842
rect 3284 842 3330 854
rect 3284 782 3290 842
rect 3324 782 3330 842
rect 3284 770 3330 782
rect 3372 842 3418 854
rect 3372 782 3378 842
rect 3412 782 3418 842
rect 3372 770 3418 782
rect 3495 842 3541 854
rect 3154 694 3200 706
rect 1405 614 1415 666
rect 1467 614 1477 666
rect 1405 608 1477 614
rect 1580 615 1590 667
rect 1642 615 1652 667
rect 2854 665 2888 694
rect 3072 665 3106 694
rect 3290 665 3324 770
rect 3495 706 3501 842
rect 3535 706 3541 842
rect 3495 694 3541 706
rect 3583 842 3629 854
rect 3583 706 3589 842
rect 3623 706 3629 842
rect 3583 694 3629 706
rect 3670 666 3704 1319
rect 3763 1224 3773 1278
rect 3825 1259 3835 1278
rect 3825 1225 4029 1259
rect 3825 1224 3835 1225
rect 3670 665 3860 666
rect 2854 631 3860 665
rect 1580 609 1652 615
rect 0 524 1424 558
rect 1458 524 3719 558
rect 340 471 350 524
rect 402 471 412 524
rect 488 496 522 524
rect 482 471 528 496
rect 482 437 488 471
rect 522 437 528 471
rect 482 412 528 437
rect 570 471 616 496
rect 570 437 576 471
rect 610 437 616 471
rect 570 412 616 437
rect 772 364 806 524
rect 846 496 880 524
rect 1022 496 1056 524
rect 1895 496 1929 524
rect 2256 496 2290 524
rect 2432 496 2466 524
rect 2762 496 2796 524
rect 3131 496 3165 524
rect 3307 496 3341 524
rect 3549 496 3583 524
rect 840 471 886 496
rect 840 437 846 471
rect 880 437 886 471
rect 840 412 886 437
rect 928 471 974 496
rect 928 437 934 471
rect 968 437 974 471
rect 928 412 974 437
rect 1016 471 1062 496
rect 1016 437 1022 471
rect 1056 437 1062 471
rect 1016 412 1062 437
rect 1418 484 1464 496
rect 1418 424 1424 484
rect 1458 424 1464 484
rect 1418 412 1464 424
rect 1506 484 1552 496
rect 1506 424 1512 484
rect 1546 424 1552 484
rect 1506 412 1552 424
rect 1594 484 1640 496
rect 1594 424 1600 484
rect 1634 424 1640 484
rect 1594 412 1640 424
rect 1889 471 1935 496
rect 1889 437 1895 471
rect 1929 437 1935 471
rect 1889 412 1935 437
rect 1977 471 2023 496
rect 1977 437 1983 471
rect 2017 437 2023 471
rect 1977 412 2023 437
rect 2250 471 2296 496
rect 2250 437 2256 471
rect 2290 437 2296 471
rect 2250 412 2296 437
rect 2338 471 2384 496
rect 2338 437 2344 471
rect 2378 437 2384 471
rect 2338 412 2384 437
rect 2426 471 2472 496
rect 2426 437 2432 471
rect 2466 437 2472 471
rect 2426 412 2472 437
rect 2514 471 2560 496
rect 2514 437 2520 471
rect 2554 437 2560 471
rect 2514 412 2560 437
rect 2756 471 2802 496
rect 2756 437 2762 471
rect 2796 437 2802 471
rect 2756 412 2802 437
rect 2844 471 2890 496
rect 2844 437 2850 471
rect 2884 437 2890 471
rect 2844 412 2890 437
rect 3125 471 3171 496
rect 3125 437 3131 471
rect 3165 437 3171 471
rect 3125 412 3171 437
rect 3213 471 3259 496
rect 3213 437 3219 471
rect 3253 437 3259 471
rect 3213 412 3259 437
rect 3301 471 3347 496
rect 3301 437 3307 471
rect 3341 437 3347 471
rect 3301 412 3347 437
rect 3543 471 3589 496
rect 3543 437 3549 471
rect 3583 437 3589 471
rect 3543 412 3589 437
rect 3631 471 3677 496
rect 3631 437 3637 471
rect 3671 437 3677 471
rect 3631 412 3677 437
rect 846 364 904 370
rect 772 330 858 364
rect 892 330 904 364
rect 846 324 904 330
rect 318 306 328 316
rect 0 272 328 306
rect 318 264 328 272
rect 380 306 390 316
rect 477 306 535 312
rect 380 272 489 306
rect 523 272 535 306
rect 380 264 390 272
rect 477 266 535 272
rect 564 306 622 312
rect 934 306 968 412
rect 1677 371 1687 396
rect 1500 365 1687 371
rect 1070 331 1512 365
rect 1546 344 1687 365
rect 1739 344 1749 396
rect 2146 350 2156 402
rect 2208 384 2218 402
rect 2344 384 2378 412
rect 2520 384 2554 412
rect 2208 365 2314 384
rect 2208 350 2268 365
rect 1546 337 1749 344
rect 1546 331 1558 337
rect 1070 306 1104 331
rect 1500 325 1558 331
rect 2256 331 2268 350
rect 2302 331 2314 365
rect 2344 350 2554 384
rect 3131 364 3189 370
rect 2256 325 2314 331
rect 1884 306 1942 312
rect 564 272 576 306
rect 610 272 738 306
rect 934 272 1104 306
rect 1707 284 1896 306
rect 1596 283 1896 284
rect 564 266 622 272
rect 704 219 738 272
rect 846 219 904 225
rect 704 185 858 219
rect 892 185 904 219
rect 846 179 904 185
rect 1021 147 1055 272
rect 1462 271 1508 283
rect 1462 211 1468 271
rect 1502 211 1508 271
rect 1462 199 1508 211
rect 1550 272 1896 283
rect 1930 272 1942 306
rect 1550 271 1735 272
rect 1550 211 1556 271
rect 1590 250 1735 271
rect 1884 266 1942 272
rect 1971 306 2029 312
rect 2520 306 2554 350
rect 3083 330 3143 364
rect 3177 330 3189 364
rect 3131 324 3189 330
rect 2751 306 2809 312
rect 1971 272 1983 306
rect 2017 294 2065 306
rect 2376 294 2434 300
rect 2017 272 2388 294
rect 1971 266 2388 272
rect 2029 260 2388 266
rect 2422 260 2434 294
rect 2376 254 2434 260
rect 2520 272 2763 306
rect 2797 272 2809 306
rect 1590 211 1596 250
rect 1550 199 1596 211
rect 2146 170 2156 222
rect 2208 213 2218 222
rect 2376 219 2434 225
rect 2376 213 2388 219
rect 2208 185 2388 213
rect 2422 185 2434 219
rect 2208 179 2434 185
rect 2208 170 2218 179
rect 2520 147 2554 272
rect 2751 266 2809 272
rect 2838 306 2896 312
rect 3219 306 3253 412
rect 3719 350 3736 402
rect 3788 350 3798 402
rect 3538 306 3596 312
rect 2838 272 2850 306
rect 2884 272 2997 306
rect 3219 272 3550 306
rect 3584 272 3596 306
rect 2838 266 2896 272
rect 2932 271 2997 272
rect 2633 219 2691 225
rect 2963 219 2997 271
rect 3131 219 3189 225
rect 2633 185 2645 219
rect 2679 185 3143 219
rect 3177 185 3189 219
rect 2633 179 2691 185
rect 482 122 528 147
rect 482 88 488 122
rect 522 88 528 122
rect 482 63 528 88
rect 570 122 616 147
rect 570 88 576 122
rect 610 88 616 122
rect 570 63 616 88
rect 840 122 886 147
rect 840 88 846 122
rect 880 88 886 122
rect 840 63 886 88
rect 928 122 974 147
rect 928 88 934 122
rect 968 88 974 122
rect 928 63 974 88
rect 1016 122 1062 147
rect 1016 88 1022 122
rect 1056 88 1062 122
rect 1016 63 1062 88
rect 1889 122 1935 147
rect 1889 88 1895 122
rect 1929 88 1935 122
rect 1889 63 1935 88
rect 1977 122 2023 147
rect 1977 88 1983 122
rect 2017 88 2023 122
rect 1977 63 2023 88
rect 2250 122 2296 147
rect 2250 88 2256 122
rect 2290 88 2296 122
rect 2250 63 2296 88
rect 2338 122 2384 147
rect 2338 88 2344 122
rect 2378 88 2384 122
rect 2338 63 2384 88
rect 2426 122 2472 147
rect 2426 88 2432 122
rect 2466 88 2472 122
rect 2426 63 2472 88
rect 2514 122 2560 147
rect 2514 88 2520 122
rect 2554 88 2560 122
rect 2514 63 2560 88
rect 2756 122 2802 147
rect 2756 88 2762 122
rect 2796 88 2802 122
rect 2756 63 2802 88
rect 2844 122 2890 147
rect 2844 88 2850 122
rect 2884 88 2890 122
rect 2844 63 2890 88
rect 2963 126 2997 185
rect 3131 179 3189 185
rect 3307 147 3341 272
rect 3538 266 3596 272
rect 3625 306 3683 312
rect 3719 306 3753 350
rect 3625 272 3637 306
rect 3671 272 3753 306
rect 3625 266 3683 272
rect 2963 73 2973 126
rect 3025 73 3035 126
rect 3125 122 3171 147
rect 3125 88 3131 122
rect 3165 88 3171 122
rect 3125 63 3171 88
rect 3213 122 3259 147
rect 3213 88 3219 122
rect 3253 88 3259 122
rect 3213 63 3259 88
rect 3301 122 3347 147
rect 3301 88 3307 122
rect 3341 88 3347 122
rect 3301 63 3347 88
rect 3543 122 3589 147
rect 3543 88 3549 122
rect 3583 88 3589 122
rect 3543 63 3589 88
rect 3631 122 3677 147
rect 3631 88 3637 122
rect 3671 88 3677 122
rect 3631 63 3677 88
rect 488 34 522 63
rect 846 34 880 63
rect 1895 34 1929 63
rect 2256 34 2290 63
rect 2762 34 2796 63
rect 3131 34 3165 63
rect 3549 34 3583 63
rect 3826 34 3860 631
rect 3914 491 4029 525
rect 3914 315 3948 491
rect 3893 263 3903 315
rect 3955 263 3965 315
rect 0 0 3860 34
<< via1 >>
rect 2477 2425 2529 2477
rect 2477 1959 2530 2011
rect 350 1789 402 1842
rect 350 1203 402 1256
rect 83 983 135 1035
rect 1415 648 1467 666
rect 1415 614 1424 648
rect 1424 614 1458 648
rect 1458 614 1467 648
rect 1590 649 1642 667
rect 1590 615 1600 649
rect 1600 615 1634 649
rect 1634 615 1642 649
rect 3773 1224 3825 1278
rect 350 471 402 524
rect 328 264 380 316
rect 1687 344 1739 396
rect 2156 350 2208 402
rect 2156 170 2208 222
rect 3736 350 3788 402
rect 2973 73 3025 126
rect 3903 263 3955 315
<< metal2 >>
rect 2477 2477 2529 2624
rect 2477 2415 2529 2425
rect 3346 2297 3398 2624
rect 1424 2263 3398 2297
rect 350 1842 402 1852
rect 350 1256 402 1789
rect 83 1035 135 1045
rect 83 973 135 983
rect 93 213 127 973
rect 350 524 402 1203
rect 1424 676 1458 2263
rect 3936 2188 3988 2624
rect 1600 2154 3988 2188
rect 1600 677 1634 2154
rect 2477 2011 2530 2021
rect 2530 1959 3912 1983
rect 2477 1949 3912 1959
rect 3773 1278 3825 1288
rect 3773 1214 3825 1224
rect 1415 666 1467 676
rect 1415 604 1467 614
rect 1590 667 1642 677
rect 1590 605 1642 615
rect 3782 507 3816 1214
rect 350 461 402 471
rect 1739 473 3816 507
rect 1739 406 1773 473
rect 3878 412 3912 1949
rect 1687 396 1773 406
rect 1739 344 1773 396
rect 1687 334 1773 344
rect 2156 402 2208 412
rect 3736 402 3912 412
rect 2208 350 3736 384
rect 3788 378 3912 402
rect 2156 340 2208 350
rect 3736 340 3788 350
rect 328 316 380 326
rect 3903 315 3955 325
rect 380 272 3903 306
rect 328 254 380 264
rect 3903 253 3955 263
rect 2156 222 2208 232
rect 93 179 2156 213
rect 2156 160 2208 170
rect 2973 126 3025 136
rect 2973 0 3025 73
<< labels >>
rlabel metal1 0 1842 34 1876 0 VDD
rlabel metal1 0 1318 34 1352 0 VSS
rlabel metal1 0 1255 34 1290 0 VDD
rlabel metal1 0 732 34 766 0 VSS
rlabel metal1 0 524 34 558 0 VDD
rlabel metal1 0 0 34 34 0 VSS
rlabel metal1 0 1590 34 1624 0 clk
rlabel metal1 0 1004 34 1038 0 cs
rlabel metal1 0 272 34 306 0 WREN
rlabel metal2 2477 2572 2529 2624 0 WLEN
rlabel metal2 3346 2572 3398 2624 0 DBL
rlabel metal2 3936 2572 3988 2624 0 DBL_
rlabel metal1 3995 1225 4029 1259 0 PCHG
rlabel metal2 2973 0 3025 53 0 SAEN
<< end >>
