.title sram_gen
.subckt bit_cell VDD VSS WL BL BL_
X0 Q Q_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X1 Q_ Q VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X2 Q Q_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 Q_ Q VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 Q WL BL VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
X5 Q_ WL BL_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
.ends bit_cell

.subckt dmy_cell VDD VSS WL BL BL_
X0 Q VSS VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X1 Q_ VDD VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X2 Q VSS VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 Q_ VDD VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 Q WL BL VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
X5 Q_ WL BL_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
.ends dmy_cell

.subckt in_reg VDD VSS clk D Q
X0 net3 clk VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X8 net3 clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 net4 net2 net5 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X10 Din net2 net1 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 net55 Q VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X13 net55 Q VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 net2 net3 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X11 net2 net3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X5 Din net3 net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X15 net4 net3 net5 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 Q net5 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X9 Q net5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X6 net11 net4 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X12 net11 net4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X7 net4 net1 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X14 net4 net1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X16 net11 net2 net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X17 net11 net3 net1 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X18 net55 net3 net5 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X19 net55 net2 net5 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X20 D_ D VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X21 D_ D VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X22 Din D_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X23 Din D_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
.ends in_reg

.subckt se_cell VDD VSS SAEN BL BL_ SB
X0 net1 SAEN VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.84
X1 diff1 BL_ net1 net1 sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X2 diff2 BL net1 net1 sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X3 diff1 diff1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 diff2 diff1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X5 diff2_ diff2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X6 diff2_ diff2 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=2
X7 SB_ diff2_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X8 SB_ diff2_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=2
X9 SB_w Q_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X10 Q_ SB_w VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.80
X11 SB_w Q_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X12 Q_ SB_w VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X13 SB_w SAEN SB_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
X14 Q_ SAEN diff2_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.60
X15 SB SB_w VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X16 SB SB_w VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
.ends se_cell

.subckt not VDD VSS A B
X0 B A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 B A VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends not

.subckt notdel VDD VSS A B
X0 B A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.84
X1 B A VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends notdel

.subckt nand2 VDD VSS A B Y
X0 Y A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 Y B VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 Y B net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X3 net1 A VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends nand2

.subckt nand3 VDD VSS A B C Y
X0 Y A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 Y B VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 Y C VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 Y A net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X4 net1 B net2 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X5 net2 C VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends nand3

.subckt nand4 VDD VSS A B C D Y
X0 Y A VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 Y B VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 Y C VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 Y D VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 Y D net1 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X5 net1 B net2 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X6 net2 C net3 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X7 net3 A VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
.ends nand4

.subckt dec_2to4 VDD VSS A1 A0 Y0 Y1 Y2 Y3
X0 VDD VSS A1 A_1 not
X1 VDD VSS A0 A_0 not
X2 VDD VSS A_1 A_0 Y0_ nand2
X3 VDD VSS A_1 A0 Y1_ nand2
X4 VDD VSS A1 A_0 Y2_ nand2
X5 VDD VSS A1 A0 Y3_ nand2
X6 VDD VSS Y0_ Y0 not
X7 VDD VSS Y1_ Y1 not
X8 VDD VSS Y2_ Y2 not
X9 VDD VSS Y3_ Y3 not
.ends dec_2to4

.subckt dec_3to6 VDD VSS A2 A1 A0 Y0 Y1 Y2 Y3 Y4 Y5
X0 VDD VSS A2 Y4 not
X1 VDD VSS Y4 Y5 not
X2 VDD VSS A1 A0 Y0 Y1 Y2 Y3 dec_2to4
.ends dec_3to6

.subckt row_dec128 VDD VSS A0 A1 A2 A3 A4 A5 A6 DC0 DC1 DC2 DC3 DC4 DC5 DC6 DC7 DC8 DC9 DC10 DC11 DC12 DC13 DC14 DC15 DC16 DC17 DC18 DC19 DC20 DC21 DC22 DC23 DC24 DC25 DC26 DC27 DC28 DC29 DC30 DC31 DC32 DC33 DC34 DC35 DC36 DC37 DC38 DC39 DC40 DC41 DC42 DC43 DC44 DC45 DC46 DC47 DC48 DC49 DC50 DC51 DC52 DC53 DC54 DC55 DC56 DC57 DC58 DC59 DC60 DC61 DC62 DC63 DC64 DC65 DC66 DC67 DC68 DC69 DC70 DC71 DC72 DC73 DC74 DC75 DC76 DC77 DC78 DC79 DC80 DC81 DC82 DC83 DC84 DC85 DC86 DC87 DC88 DC89 DC90 DC91 DC92 DC93 DC94 DC95 DC96 DC97 DC98 DC99 DC100 DC101 DC102 DC103 DC104 DC105 DC106 DC107 DC108 DC109 DC110 DC111 DC112 DC113 DC114 DC115 DC116 DC117 DC118 DC119 DC120 DC121 DC122 DC123 DC124 DC125 DC126 DC127
X0 VDD VSS A1 A0 Y0 Y1 Y2 Y3 dec_2to4
X1 VDD VSS A3 A2 Y4 Y5 Y6 Y7 dec_2to4
X2 VDD VSS A6 A5 A4 Y8 Y9 Y10 Y11 Y12 Y13 dec_3to6
X3 VDD VSS Y0 Y4 Y8 Y12 DC_0 nand4
X4 VDD VSS Y1 Y4 Y8 Y12 DC_1 nand4
X5 VDD VSS Y2 Y4 Y8 Y12 DC_2 nand4
X6 VDD VSS Y3 Y4 Y8 Y12 DC_3 nand4
X7 VDD VSS Y0 Y5 Y8 Y12 DC_4 nand4
X8 VDD VSS Y1 Y5 Y8 Y12 DC_5 nand4
X9 VDD VSS Y2 Y5 Y8 Y12 DC_6 nand4
X10 VDD VSS Y3 Y5 Y8 Y12 DC_7 nand4
X11 VDD VSS Y0 Y6 Y8 Y12 DC_8 nand4
X12 VDD VSS Y1 Y6 Y8 Y12 DC_9 nand4
X13 VDD VSS Y2 Y6 Y8 Y12 DC_10 nand4
X14 VDD VSS Y3 Y6 Y8 Y12 DC_11 nand4
X15 VDD VSS Y0 Y7 Y8 Y12 DC_12 nand4
X16 VDD VSS Y1 Y7 Y8 Y12 DC_13 nand4
X17 VDD VSS Y2 Y7 Y8 Y12 DC_14 nand4
X18 VDD VSS Y3 Y7 Y8 Y12 DC_15 nand4
X19 VDD VSS Y0 Y4 Y9 Y12 DC_16 nand4
X20 VDD VSS Y1 Y4 Y9 Y12 DC_17 nand4
X21 VDD VSS Y2 Y4 Y9 Y12 DC_18 nand4
X22 VDD VSS Y3 Y4 Y9 Y12 DC_19 nand4
X23 VDD VSS Y0 Y5 Y9 Y12 DC_20 nand4
X24 VDD VSS Y1 Y5 Y9 Y12 DC_21 nand4
X25 VDD VSS Y2 Y5 Y9 Y12 DC_22 nand4
X26 VDD VSS Y3 Y5 Y9 Y12 DC_23 nand4
X27 VDD VSS Y0 Y6 Y9 Y12 DC_24 nand4
X28 VDD VSS Y1 Y6 Y9 Y12 DC_25 nand4
X29 VDD VSS Y2 Y6 Y9 Y12 DC_26 nand4
X30 VDD VSS Y3 Y6 Y9 Y12 DC_27 nand4
X31 VDD VSS Y0 Y7 Y9 Y12 DC_28 nand4
X32 VDD VSS Y1 Y7 Y9 Y12 DC_29 nand4
X33 VDD VSS Y2 Y7 Y9 Y12 DC_30 nand4
X34 VDD VSS Y3 Y7 Y9 Y12 DC_31 nand4
X35 VDD VSS Y0 Y4 Y10 Y12 DC_32 nand4
X36 VDD VSS Y1 Y4 Y10 Y12 DC_33 nand4
X37 VDD VSS Y2 Y4 Y10 Y12 DC_34 nand4
X38 VDD VSS Y3 Y4 Y10 Y12 DC_35 nand4
X39 VDD VSS Y0 Y5 Y10 Y12 DC_36 nand4
X40 VDD VSS Y1 Y5 Y10 Y12 DC_37 nand4
X41 VDD VSS Y2 Y5 Y10 Y12 DC_38 nand4
X42 VDD VSS Y3 Y5 Y10 Y12 DC_39 nand4
X43 VDD VSS Y0 Y6 Y10 Y12 DC_40 nand4
X44 VDD VSS Y1 Y6 Y10 Y12 DC_41 nand4
X45 VDD VSS Y2 Y6 Y10 Y12 DC_42 nand4
X46 VDD VSS Y3 Y6 Y10 Y12 DC_43 nand4
X47 VDD VSS Y0 Y7 Y10 Y12 DC_44 nand4
X48 VDD VSS Y1 Y7 Y10 Y12 DC_45 nand4
X49 VDD VSS Y2 Y7 Y10 Y12 DC_46 nand4
X50 VDD VSS Y3 Y7 Y10 Y12 DC_47 nand4
X51 VDD VSS Y0 Y4 Y11 Y12 DC_48 nand4
X52 VDD VSS Y1 Y4 Y11 Y12 DC_49 nand4
X53 VDD VSS Y2 Y4 Y11 Y12 DC_50 nand4
X54 VDD VSS Y3 Y4 Y11 Y12 DC_51 nand4
X55 VDD VSS Y0 Y5 Y11 Y12 DC_52 nand4
X56 VDD VSS Y1 Y5 Y11 Y12 DC_53 nand4
X57 VDD VSS Y2 Y5 Y11 Y12 DC_54 nand4
X58 VDD VSS Y3 Y5 Y11 Y12 DC_55 nand4
X59 VDD VSS Y0 Y6 Y11 Y12 DC_56 nand4
X60 VDD VSS Y1 Y6 Y11 Y12 DC_57 nand4
X61 VDD VSS Y2 Y6 Y11 Y12 DC_58 nand4
X62 VDD VSS Y3 Y6 Y11 Y12 DC_59 nand4
X63 VDD VSS Y0 Y7 Y11 Y12 DC_60 nand4
X64 VDD VSS Y1 Y7 Y11 Y12 DC_61 nand4
X65 VDD VSS Y2 Y7 Y11 Y12 DC_62 nand4
X66 VDD VSS Y3 Y7 Y11 Y12 DC_63 nand4
X67 VDD VSS Y0 Y4 Y8 Y13 DC_64 nand4
X68 VDD VSS Y1 Y4 Y8 Y13 DC_65 nand4
X69 VDD VSS Y2 Y4 Y8 Y13 DC_66 nand4
X70 VDD VSS Y3 Y4 Y8 Y13 DC_67 nand4
X71 VDD VSS Y0 Y5 Y8 Y13 DC_68 nand4
X72 VDD VSS Y1 Y5 Y8 Y13 DC_69 nand4
X73 VDD VSS Y2 Y5 Y8 Y13 DC_70 nand4
X74 VDD VSS Y3 Y5 Y8 Y13 DC_71 nand4
X75 VDD VSS Y0 Y6 Y8 Y13 DC_72 nand4
X76 VDD VSS Y1 Y6 Y8 Y13 DC_73 nand4
X77 VDD VSS Y2 Y6 Y8 Y13 DC_74 nand4
X78 VDD VSS Y3 Y6 Y8 Y13 DC_75 nand4
X79 VDD VSS Y0 Y7 Y8 Y13 DC_76 nand4
X80 VDD VSS Y1 Y7 Y8 Y13 DC_77 nand4
X81 VDD VSS Y2 Y7 Y8 Y13 DC_78 nand4
X82 VDD VSS Y3 Y7 Y8 Y13 DC_79 nand4
X83 VDD VSS Y0 Y4 Y9 Y13 DC_80 nand4
X84 VDD VSS Y1 Y4 Y9 Y13 DC_81 nand4
X85 VDD VSS Y2 Y4 Y9 Y13 DC_82 nand4
X86 VDD VSS Y3 Y4 Y9 Y13 DC_83 nand4
X87 VDD VSS Y0 Y5 Y9 Y13 DC_84 nand4
X88 VDD VSS Y1 Y5 Y9 Y13 DC_85 nand4
X89 VDD VSS Y2 Y5 Y9 Y13 DC_86 nand4
X90 VDD VSS Y3 Y5 Y9 Y13 DC_87 nand4
X91 VDD VSS Y0 Y6 Y9 Y13 DC_88 nand4
X92 VDD VSS Y1 Y6 Y9 Y13 DC_89 nand4
X93 VDD VSS Y2 Y6 Y9 Y13 DC_90 nand4
X94 VDD VSS Y3 Y6 Y9 Y13 DC_91 nand4
X95 VDD VSS Y0 Y7 Y9 Y13 DC_92 nand4
X96 VDD VSS Y1 Y7 Y9 Y13 DC_93 nand4
X97 VDD VSS Y2 Y7 Y9 Y13 DC_94 nand4
X98 VDD VSS Y3 Y7 Y9 Y13 DC_95 nand4
X99 VDD VSS Y0 Y4 Y10 Y13 DC_96 nand4
X100 VDD VSS Y1 Y4 Y10 Y13 DC_97 nand4
X101 VDD VSS Y2 Y4 Y10 Y13 DC_98 nand4
X102 VDD VSS Y3 Y4 Y10 Y13 DC_99 nand4
X103 VDD VSS Y0 Y5 Y10 Y13 DC_100 nand4
X104 VDD VSS Y1 Y5 Y10 Y13 DC_101 nand4
X105 VDD VSS Y2 Y5 Y10 Y13 DC_102 nand4
X106 VDD VSS Y3 Y5 Y10 Y13 DC_103 nand4
X107 VDD VSS Y0 Y6 Y10 Y13 DC_104 nand4
X108 VDD VSS Y1 Y6 Y10 Y13 DC_105 nand4
X109 VDD VSS Y2 Y6 Y10 Y13 DC_106 nand4
X110 VDD VSS Y3 Y6 Y10 Y13 DC_107 nand4
X111 VDD VSS Y0 Y7 Y10 Y13 DC_108 nand4
X112 VDD VSS Y1 Y7 Y10 Y13 DC_109 nand4
X113 VDD VSS Y2 Y7 Y10 Y13 DC_110 nand4
X114 VDD VSS Y3 Y7 Y10 Y13 DC_111 nand4
X115 VDD VSS Y0 Y4 Y11 Y13 DC_112 nand4
X116 VDD VSS Y1 Y4 Y11 Y13 DC_113 nand4
X117 VDD VSS Y2 Y4 Y11 Y13 DC_114 nand4
X118 VDD VSS Y3 Y4 Y11 Y13 DC_115 nand4
X119 VDD VSS Y0 Y5 Y11 Y13 DC_116 nand4
X120 VDD VSS Y1 Y5 Y11 Y13 DC_117 nand4
X121 VDD VSS Y2 Y5 Y11 Y13 DC_118 nand4
X122 VDD VSS Y3 Y5 Y11 Y13 DC_119 nand4
X123 VDD VSS Y0 Y6 Y11 Y13 DC_120 nand4
X124 VDD VSS Y1 Y6 Y11 Y13 DC_121 nand4
X125 VDD VSS Y2 Y6 Y11 Y13 DC_122 nand4
X126 VDD VSS Y3 Y6 Y11 Y13 DC_123 nand4
X127 VDD VSS Y0 Y7 Y11 Y13 DC_124 nand4
X128 VDD VSS Y1 Y7 Y11 Y13 DC_125 nand4
X129 VDD VSS Y2 Y7 Y11 Y13 DC_126 nand4
X130 VDD VSS Y3 Y7 Y11 Y13 DC_127 nand4
X131 VDD VSS DC_0 DC0 not
X132 VDD VSS DC_1 DC1 not
X133 VDD VSS DC_2 DC2 not
X134 VDD VSS DC_3 DC3 not
X135 VDD VSS DC_4 DC4 not
X136 VDD VSS DC_5 DC5 not
X137 VDD VSS DC_6 DC6 not
X138 VDD VSS DC_7 DC7 not
X139 VDD VSS DC_8 DC8 not
X140 VDD VSS DC_9 DC9 not
X141 VDD VSS DC_10 DC10 not
X142 VDD VSS DC_11 DC11 not
X143 VDD VSS DC_12 DC12 not
X144 VDD VSS DC_13 DC13 not
X145 VDD VSS DC_14 DC14 not
X146 VDD VSS DC_15 DC15 not
X147 VDD VSS DC_16 DC16 not
X148 VDD VSS DC_17 DC17 not
X149 VDD VSS DC_18 DC18 not
X150 VDD VSS DC_19 DC19 not
X151 VDD VSS DC_20 DC20 not
X152 VDD VSS DC_21 DC21 not
X153 VDD VSS DC_22 DC22 not
X154 VDD VSS DC_23 DC23 not
X155 VDD VSS DC_24 DC24 not
X156 VDD VSS DC_25 DC25 not
X157 VDD VSS DC_26 DC26 not
X158 VDD VSS DC_27 DC27 not
X159 VDD VSS DC_28 DC28 not
X160 VDD VSS DC_29 DC29 not
X161 VDD VSS DC_30 DC30 not
X162 VDD VSS DC_31 DC31 not
X163 VDD VSS DC_32 DC32 not
X164 VDD VSS DC_33 DC33 not
X165 VDD VSS DC_34 DC34 not
X166 VDD VSS DC_35 DC35 not
X167 VDD VSS DC_36 DC36 not
X168 VDD VSS DC_37 DC37 not
X169 VDD VSS DC_38 DC38 not
X170 VDD VSS DC_39 DC39 not
X171 VDD VSS DC_40 DC40 not
X172 VDD VSS DC_41 DC41 not
X173 VDD VSS DC_42 DC42 not
X174 VDD VSS DC_43 DC43 not
X175 VDD VSS DC_44 DC44 not
X176 VDD VSS DC_45 DC45 not
X177 VDD VSS DC_46 DC46 not
X178 VDD VSS DC_47 DC47 not
X179 VDD VSS DC_48 DC48 not
X180 VDD VSS DC_49 DC49 not
X181 VDD VSS DC_50 DC50 not
X182 VDD VSS DC_51 DC51 not
X183 VDD VSS DC_52 DC52 not
X184 VDD VSS DC_53 DC53 not
X185 VDD VSS DC_54 DC54 not
X186 VDD VSS DC_55 DC55 not
X187 VDD VSS DC_56 DC56 not
X188 VDD VSS DC_57 DC57 not
X189 VDD VSS DC_58 DC58 not
X190 VDD VSS DC_59 DC59 not
X191 VDD VSS DC_60 DC60 not
X192 VDD VSS DC_61 DC61 not
X193 VDD VSS DC_62 DC62 not
X194 VDD VSS DC_63 DC63 not
X195 VDD VSS DC_64 DC64 not
X196 VDD VSS DC_65 DC65 not
X197 VDD VSS DC_66 DC66 not
X198 VDD VSS DC_67 DC67 not
X199 VDD VSS DC_68 DC68 not
X200 VDD VSS DC_69 DC69 not
X201 VDD VSS DC_70 DC70 not
X202 VDD VSS DC_71 DC71 not
X203 VDD VSS DC_72 DC72 not
X204 VDD VSS DC_73 DC73 not
X205 VDD VSS DC_74 DC74 not
X206 VDD VSS DC_75 DC75 not
X207 VDD VSS DC_76 DC76 not
X208 VDD VSS DC_77 DC77 not
X209 VDD VSS DC_78 DC78 not
X210 VDD VSS DC_79 DC79 not
X211 VDD VSS DC_80 DC80 not
X212 VDD VSS DC_81 DC81 not
X213 VDD VSS DC_82 DC82 not
X214 VDD VSS DC_83 DC83 not
X215 VDD VSS DC_84 DC84 not
X216 VDD VSS DC_85 DC85 not
X217 VDD VSS DC_86 DC86 not
X218 VDD VSS DC_87 DC87 not
X219 VDD VSS DC_88 DC88 not
X220 VDD VSS DC_89 DC89 not
X221 VDD VSS DC_90 DC90 not
X222 VDD VSS DC_91 DC91 not
X223 VDD VSS DC_92 DC92 not
X224 VDD VSS DC_93 DC93 not
X225 VDD VSS DC_94 DC94 not
X226 VDD VSS DC_95 DC95 not
X227 VDD VSS DC_96 DC96 not
X228 VDD VSS DC_97 DC97 not
X229 VDD VSS DC_98 DC98 not
X230 VDD VSS DC_99 DC99 not
X231 VDD VSS DC_100 DC100 not
X232 VDD VSS DC_101 DC101 not
X233 VDD VSS DC_102 DC102 not
X234 VDD VSS DC_103 DC103 not
X235 VDD VSS DC_104 DC104 not
X236 VDD VSS DC_105 DC105 not
X237 VDD VSS DC_106 DC106 not
X238 VDD VSS DC_107 DC107 not
X239 VDD VSS DC_108 DC108 not
X240 VDD VSS DC_109 DC109 not
X241 VDD VSS DC_110 DC110 not
X242 VDD VSS DC_111 DC111 not
X243 VDD VSS DC_112 DC112 not
X244 VDD VSS DC_113 DC113 not
X245 VDD VSS DC_114 DC114 not
X246 VDD VSS DC_115 DC115 not
X247 VDD VSS DC_116 DC116 not
X248 VDD VSS DC_117 DC117 not
X249 VDD VSS DC_118 DC118 not
X250 VDD VSS DC_119 DC119 not
X251 VDD VSS DC_120 DC120 not
X252 VDD VSS DC_121 DC121 not
X253 VDD VSS DC_122 DC122 not
X254 VDD VSS DC_123 DC123 not
X255 VDD VSS DC_124 DC124 not
X256 VDD VSS DC_125 DC125 not
X257 VDD VSS DC_126 DC126 not
X258 VDD VSS DC_127 DC127 not
.ends row_dec128

.subckt row_driver VDD VSS WLEN A B
X0 VDD VSS A WLEN net1 nand2
X1 B net1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X2 B net1 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
.ends row_driver

.subckt rd_arr_128 VDD VSS WLEN DC0 DC1 DC2 DC3 DC4 DC5 DC6 DC7 DC8 DC9 DC10 DC11 DC12 DC13 DC14 DC15 DC16 DC17 DC18 DC19 DC20 DC21 DC22 DC23 DC24 DC25 DC26 DC27 DC28 DC29 DC30 DC31 DC32 DC33 DC34 DC35 DC36 DC37 DC38 DC39 DC40 DC41 DC42 DC43 DC44 DC45 DC46 DC47 DC48 DC49 DC50 DC51 DC52 DC53 DC54 DC55 DC56 DC57 DC58 DC59 DC60 DC61 DC62 DC63 DC64 DC65 DC66 DC67 DC68 DC69 DC70 DC71 DC72 DC73 DC74 DC75 DC76 DC77 DC78 DC79 DC80 DC81 DC82 DC83 DC84 DC85 DC86 DC87 DC88 DC89 DC90 DC91 DC92 DC93 DC94 DC95 DC96 DC97 DC98 DC99 DC100 DC101 DC102 DC103 DC104 DC105 DC106 DC107 DC108 DC109 DC110 DC111 DC112 DC113 DC114 DC115 DC116 DC117 DC118 DC119 DC120 DC121 DC122 DC123 DC124 DC125 DC126 DC127 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 WL32 WL33 WL34 WL35 WL36 WL37 WL38 WL39 WL40 WL41 WL42 WL43 WL44 WL45 WL46 WL47 WL48 WL49 WL50 WL51 WL52 WL53 WL54 WL55 WL56 WL57 WL58 WL59 WL60 WL61 WL62 WL63 WL64 WL65 WL66 WL67 WL68 WL69 WL70 WL71 WL72 WL73 WL74 WL75 WL76 WL77 WL78 WL79 WL80 WL81 WL82 WL83 WL84 WL85 WL86 WL87 WL88 WL89 WL90 WL91 WL92 WL93 WL94 WL95 WL96 WL97 WL98 WL99 WL100 WL101 WL102 WL103 WL104 WL105 WL106 WL107 WL108 WL109 WL110 WL111 WL112 WL113 WL114 WL115 WL116 WL117 WL118 WL119 WL120 WL121 WL122 WL123 WL124 WL125 WL126 WL127
X0 VDD VSS WLEN DC0 WL0 row_driver
X1 VDD VSS WLEN DC1 WL1 row_driver
X2 VDD VSS WLEN DC2 WL2 row_driver
X3 VDD VSS WLEN DC3 WL3 row_driver
X4 VDD VSS WLEN DC4 WL4 row_driver
X5 VDD VSS WLEN DC5 WL5 row_driver
X6 VDD VSS WLEN DC6 WL6 row_driver
X7 VDD VSS WLEN DC7 WL7 row_driver
X8 VDD VSS WLEN DC8 WL8 row_driver
X9 VDD VSS WLEN DC9 WL9 row_driver
X10 VDD VSS WLEN DC10 WL10 row_driver
X11 VDD VSS WLEN DC11 WL11 row_driver
X12 VDD VSS WLEN DC12 WL12 row_driver
X13 VDD VSS WLEN DC13 WL13 row_driver
X14 VDD VSS WLEN DC14 WL14 row_driver
X15 VDD VSS WLEN DC15 WL15 row_driver
X16 VDD VSS WLEN DC16 WL16 row_driver
X17 VDD VSS WLEN DC17 WL17 row_driver
X18 VDD VSS WLEN DC18 WL18 row_driver
X19 VDD VSS WLEN DC19 WL19 row_driver
X20 VDD VSS WLEN DC20 WL20 row_driver
X21 VDD VSS WLEN DC21 WL21 row_driver
X22 VDD VSS WLEN DC22 WL22 row_driver
X23 VDD VSS WLEN DC23 WL23 row_driver
X24 VDD VSS WLEN DC24 WL24 row_driver
X25 VDD VSS WLEN DC25 WL25 row_driver
X26 VDD VSS WLEN DC26 WL26 row_driver
X27 VDD VSS WLEN DC27 WL27 row_driver
X28 VDD VSS WLEN DC28 WL28 row_driver
X29 VDD VSS WLEN DC29 WL29 row_driver
X30 VDD VSS WLEN DC30 WL30 row_driver
X31 VDD VSS WLEN DC31 WL31 row_driver
X32 VDD VSS WLEN DC32 WL32 row_driver
X33 VDD VSS WLEN DC33 WL33 row_driver
X34 VDD VSS WLEN DC34 WL34 row_driver
X35 VDD VSS WLEN DC35 WL35 row_driver
X36 VDD VSS WLEN DC36 WL36 row_driver
X37 VDD VSS WLEN DC37 WL37 row_driver
X38 VDD VSS WLEN DC38 WL38 row_driver
X39 VDD VSS WLEN DC39 WL39 row_driver
X40 VDD VSS WLEN DC40 WL40 row_driver
X41 VDD VSS WLEN DC41 WL41 row_driver
X42 VDD VSS WLEN DC42 WL42 row_driver
X43 VDD VSS WLEN DC43 WL43 row_driver
X44 VDD VSS WLEN DC44 WL44 row_driver
X45 VDD VSS WLEN DC45 WL45 row_driver
X46 VDD VSS WLEN DC46 WL46 row_driver
X47 VDD VSS WLEN DC47 WL47 row_driver
X48 VDD VSS WLEN DC48 WL48 row_driver
X49 VDD VSS WLEN DC49 WL49 row_driver
X50 VDD VSS WLEN DC50 WL50 row_driver
X51 VDD VSS WLEN DC51 WL51 row_driver
X52 VDD VSS WLEN DC52 WL52 row_driver
X53 VDD VSS WLEN DC53 WL53 row_driver
X54 VDD VSS WLEN DC54 WL54 row_driver
X55 VDD VSS WLEN DC55 WL55 row_driver
X56 VDD VSS WLEN DC56 WL56 row_driver
X57 VDD VSS WLEN DC57 WL57 row_driver
X58 VDD VSS WLEN DC58 WL58 row_driver
X59 VDD VSS WLEN DC59 WL59 row_driver
X60 VDD VSS WLEN DC60 WL60 row_driver
X61 VDD VSS WLEN DC61 WL61 row_driver
X62 VDD VSS WLEN DC62 WL62 row_driver
X63 VDD VSS WLEN DC63 WL63 row_driver
X64 VDD VSS WLEN DC64 WL64 row_driver
X65 VDD VSS WLEN DC65 WL65 row_driver
X66 VDD VSS WLEN DC66 WL66 row_driver
X67 VDD VSS WLEN DC67 WL67 row_driver
X68 VDD VSS WLEN DC68 WL68 row_driver
X69 VDD VSS WLEN DC69 WL69 row_driver
X70 VDD VSS WLEN DC70 WL70 row_driver
X71 VDD VSS WLEN DC71 WL71 row_driver
X72 VDD VSS WLEN DC72 WL72 row_driver
X73 VDD VSS WLEN DC73 WL73 row_driver
X74 VDD VSS WLEN DC74 WL74 row_driver
X75 VDD VSS WLEN DC75 WL75 row_driver
X76 VDD VSS WLEN DC76 WL76 row_driver
X77 VDD VSS WLEN DC77 WL77 row_driver
X78 VDD VSS WLEN DC78 WL78 row_driver
X79 VDD VSS WLEN DC79 WL79 row_driver
X80 VDD VSS WLEN DC80 WL80 row_driver
X81 VDD VSS WLEN DC81 WL81 row_driver
X82 VDD VSS WLEN DC82 WL82 row_driver
X83 VDD VSS WLEN DC83 WL83 row_driver
X84 VDD VSS WLEN DC84 WL84 row_driver
X85 VDD VSS WLEN DC85 WL85 row_driver
X86 VDD VSS WLEN DC86 WL86 row_driver
X87 VDD VSS WLEN DC87 WL87 row_driver
X88 VDD VSS WLEN DC88 WL88 row_driver
X89 VDD VSS WLEN DC89 WL89 row_driver
X90 VDD VSS WLEN DC90 WL90 row_driver
X91 VDD VSS WLEN DC91 WL91 row_driver
X92 VDD VSS WLEN DC92 WL92 row_driver
X93 VDD VSS WLEN DC93 WL93 row_driver
X94 VDD VSS WLEN DC94 WL94 row_driver
X95 VDD VSS WLEN DC95 WL95 row_driver
X96 VDD VSS WLEN DC96 WL96 row_driver
X97 VDD VSS WLEN DC97 WL97 row_driver
X98 VDD VSS WLEN DC98 WL98 row_driver
X99 VDD VSS WLEN DC99 WL99 row_driver
X100 VDD VSS WLEN DC100 WL100 row_driver
X101 VDD VSS WLEN DC101 WL101 row_driver
X102 VDD VSS WLEN DC102 WL102 row_driver
X103 VDD VSS WLEN DC103 WL103 row_driver
X104 VDD VSS WLEN DC104 WL104 row_driver
X105 VDD VSS WLEN DC105 WL105 row_driver
X106 VDD VSS WLEN DC106 WL106 row_driver
X107 VDD VSS WLEN DC107 WL107 row_driver
X108 VDD VSS WLEN DC108 WL108 row_driver
X109 VDD VSS WLEN DC109 WL109 row_driver
X110 VDD VSS WLEN DC110 WL110 row_driver
X111 VDD VSS WLEN DC111 WL111 row_driver
X112 VDD VSS WLEN DC112 WL112 row_driver
X113 VDD VSS WLEN DC113 WL113 row_driver
X114 VDD VSS WLEN DC114 WL114 row_driver
X115 VDD VSS WLEN DC115 WL115 row_driver
X116 VDD VSS WLEN DC116 WL116 row_driver
X117 VDD VSS WLEN DC117 WL117 row_driver
X118 VDD VSS WLEN DC118 WL118 row_driver
X119 VDD VSS WLEN DC119 WL119 row_driver
X120 VDD VSS WLEN DC120 WL120 row_driver
X121 VDD VSS WLEN DC121 WL121 row_driver
X122 VDD VSS WLEN DC122 WL122 row_driver
X123 VDD VSS WLEN DC123 WL123 row_driver
X124 VDD VSS WLEN DC124 WL124 row_driver
X125 VDD VSS WLEN DC125 WL125 row_driver
X126 VDD VSS WLEN DC126 WL126 row_driver
X127 VDD VSS WLEN DC127 WL127 row_driver
.ends rd_arr_128

.subckt col_dec1 VDD VSS DC0
X0 DC0 VDD VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X1 DC0 VDD VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
.ends col_dec1

.subckt dido VDD VSS PCHG WREN SEL BL BL_ DW DW_ DR DR_
X0 BL_ net6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 BL net6 BL_ VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X2 BL net6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 net6 net5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X4 net6 net5 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X5 net5 PCHG VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X6 net5 PCHG VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X7 BL_ net3 DR_ VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X8 DR net3 BL VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X9 net4 SEL VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X10 BL net2 DW VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X11 DW_ net2 BL_ VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X12 net4 SEL VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X13 net3 net4 VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X14 net3 net4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X15 VDD VSS net4 WREN net1 nand2
X16 VDD VSS net1 net2 not
.ends dido

.subckt dido_arr_64 VDD VSS PCHG WREN SEL0 SEL1 SEL2 SEL3 SEL4 SEL5 SEL6 SEL7 SEL8 SEL9 SEL10 SEL11 SEL12 SEL13 SEL14 SEL15 SEL16 SEL17 SEL18 SEL19 SEL20 SEL21 SEL22 SEL23 SEL24 SEL25 SEL26 SEL27 SEL28 SEL29 SEL30 SEL31 SEL32 SEL33 SEL34 SEL35 SEL36 SEL37 SEL38 SEL39 SEL40 SEL41 SEL42 SEL43 SEL44 SEL45 SEL46 SEL47 SEL48 SEL49 SEL50 SEL51 SEL52 SEL53 SEL54 SEL55 SEL56 SEL57 SEL58 SEL59 SEL60 SEL61 SEL62 SEL63 BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 DW0 DW_0 DW1 DW_1 DW2 DW_2 DW3 DW_3 DW4 DW_4 DW5 DW_5 DW6 DW_6 DW7 DW_7 DW8 DW_8 DW9 DW_9 DW10 DW_10 DW11 DW_11 DW12 DW_12 DW13 DW_13 DW14 DW_14 DW15 DW_15 DW16 DW_16 DW17 DW_17 DW18 DW_18 DW19 DW_19 DW20 DW_20 DW21 DW_21 DW22 DW_22 DW23 DW_23 DW24 DW_24 DW25 DW_25 DW26 DW_26 DW27 DW_27 DW28 DW_28 DW29 DW_29 DW30 DW_30 DW31 DW_31 DW32 DW_32 DW33 DW_33 DW34 DW_34 DW35 DW_35 DW36 DW_36 DW37 DW_37 DW38 DW_38 DW39 DW_39 DW40 DW_40 DW41 DW_41 DW42 DW_42 DW43 DW_43 DW44 DW_44 DW45 DW_45 DW46 DW_46 DW47 DW_47 DW48 DW_48 DW49 DW_49 DW50 DW_50 DW51 DW_51 DW52 DW_52 DW53 DW_53 DW54 DW_54 DW55 DW_55 DW56 DW_56 DW57 DW_57 DW58 DW_58 DW59 DW_59 DW60 DW_60 DW61 DW_61 DW62 DW_62 DW63 DW_63 DR0 DR_0 DR1 DR_1 DR2 DR_2 DR3 DR_3 DR4 DR_4 DR5 DR_5 DR6 DR_6 DR7 DR_7 DR8 DR_8 DR9 DR_9 DR10 DR_10 DR11 DR_11 DR12 DR_12 DR13 DR_13 DR14 DR_14 DR15 DR_15 DR16 DR_16 DR17 DR_17 DR18 DR_18 DR19 DR_19 DR20 DR_20 DR21 DR_21 DR22 DR_22 DR23 DR_23 DR24 DR_24 DR25 DR_25 DR26 DR_26 DR27 DR_27 DR28 DR_28 DR29 DR_29 DR30 DR_30 DR31 DR_31 DR32 DR_32 DR33 DR_33 DR34 DR_34 DR35 DR_35 DR36 DR_36 DR37 DR_37 DR38 DR_38 DR39 DR_39 DR40 DR_40 DR41 DR_41 DR42 DR_42 DR43 DR_43 DR44 DR_44 DR45 DR_45 DR46 DR_46 DR47 DR_47 DR48 DR_48 DR49 DR_49 DR50 DR_50 DR51 DR_51 DR52 DR_52 DR53 DR_53 DR54 DR_54 DR55 DR_55 DR56 DR_56 DR57 DR_57 DR58 DR_58 DR59 DR_59 DR60 DR_60 DR61 DR_61 DR62 DR_62 DR63 DR_63
X0 VDD VSS PCHG WREN SEL0 BL0 BL_0 DW0 DW_0 DR0 DR_0 dido
X1 VDD VSS PCHG WREN SEL1 BL1 BL_1 DW1 DW_1 DR1 DR_1 dido
X2 VDD VSS PCHG WREN SEL2 BL2 BL_2 DW2 DW_2 DR2 DR_2 dido
X3 VDD VSS PCHG WREN SEL3 BL3 BL_3 DW3 DW_3 DR3 DR_3 dido
X4 VDD VSS PCHG WREN SEL4 BL4 BL_4 DW4 DW_4 DR4 DR_4 dido
X5 VDD VSS PCHG WREN SEL5 BL5 BL_5 DW5 DW_5 DR5 DR_5 dido
X6 VDD VSS PCHG WREN SEL6 BL6 BL_6 DW6 DW_6 DR6 DR_6 dido
X7 VDD VSS PCHG WREN SEL7 BL7 BL_7 DW7 DW_7 DR7 DR_7 dido
X8 VDD VSS PCHG WREN SEL8 BL8 BL_8 DW8 DW_8 DR8 DR_8 dido
X9 VDD VSS PCHG WREN SEL9 BL9 BL_9 DW9 DW_9 DR9 DR_9 dido
X10 VDD VSS PCHG WREN SEL10 BL10 BL_10 DW10 DW_10 DR10 DR_10 dido
X11 VDD VSS PCHG WREN SEL11 BL11 BL_11 DW11 DW_11 DR11 DR_11 dido
X12 VDD VSS PCHG WREN SEL12 BL12 BL_12 DW12 DW_12 DR12 DR_12 dido
X13 VDD VSS PCHG WREN SEL13 BL13 BL_13 DW13 DW_13 DR13 DR_13 dido
X14 VDD VSS PCHG WREN SEL14 BL14 BL_14 DW14 DW_14 DR14 DR_14 dido
X15 VDD VSS PCHG WREN SEL15 BL15 BL_15 DW15 DW_15 DR15 DR_15 dido
X16 VDD VSS PCHG WREN SEL16 BL16 BL_16 DW16 DW_16 DR16 DR_16 dido
X17 VDD VSS PCHG WREN SEL17 BL17 BL_17 DW17 DW_17 DR17 DR_17 dido
X18 VDD VSS PCHG WREN SEL18 BL18 BL_18 DW18 DW_18 DR18 DR_18 dido
X19 VDD VSS PCHG WREN SEL19 BL19 BL_19 DW19 DW_19 DR19 DR_19 dido
X20 VDD VSS PCHG WREN SEL20 BL20 BL_20 DW20 DW_20 DR20 DR_20 dido
X21 VDD VSS PCHG WREN SEL21 BL21 BL_21 DW21 DW_21 DR21 DR_21 dido
X22 VDD VSS PCHG WREN SEL22 BL22 BL_22 DW22 DW_22 DR22 DR_22 dido
X23 VDD VSS PCHG WREN SEL23 BL23 BL_23 DW23 DW_23 DR23 DR_23 dido
X24 VDD VSS PCHG WREN SEL24 BL24 BL_24 DW24 DW_24 DR24 DR_24 dido
X25 VDD VSS PCHG WREN SEL25 BL25 BL_25 DW25 DW_25 DR25 DR_25 dido
X26 VDD VSS PCHG WREN SEL26 BL26 BL_26 DW26 DW_26 DR26 DR_26 dido
X27 VDD VSS PCHG WREN SEL27 BL27 BL_27 DW27 DW_27 DR27 DR_27 dido
X28 VDD VSS PCHG WREN SEL28 BL28 BL_28 DW28 DW_28 DR28 DR_28 dido
X29 VDD VSS PCHG WREN SEL29 BL29 BL_29 DW29 DW_29 DR29 DR_29 dido
X30 VDD VSS PCHG WREN SEL30 BL30 BL_30 DW30 DW_30 DR30 DR_30 dido
X31 VDD VSS PCHG WREN SEL31 BL31 BL_31 DW31 DW_31 DR31 DR_31 dido
X32 VDD VSS PCHG WREN SEL32 BL32 BL_32 DW32 DW_32 DR32 DR_32 dido
X33 VDD VSS PCHG WREN SEL33 BL33 BL_33 DW33 DW_33 DR33 DR_33 dido
X34 VDD VSS PCHG WREN SEL34 BL34 BL_34 DW34 DW_34 DR34 DR_34 dido
X35 VDD VSS PCHG WREN SEL35 BL35 BL_35 DW35 DW_35 DR35 DR_35 dido
X36 VDD VSS PCHG WREN SEL36 BL36 BL_36 DW36 DW_36 DR36 DR_36 dido
X37 VDD VSS PCHG WREN SEL37 BL37 BL_37 DW37 DW_37 DR37 DR_37 dido
X38 VDD VSS PCHG WREN SEL38 BL38 BL_38 DW38 DW_38 DR38 DR_38 dido
X39 VDD VSS PCHG WREN SEL39 BL39 BL_39 DW39 DW_39 DR39 DR_39 dido
X40 VDD VSS PCHG WREN SEL40 BL40 BL_40 DW40 DW_40 DR40 DR_40 dido
X41 VDD VSS PCHG WREN SEL41 BL41 BL_41 DW41 DW_41 DR41 DR_41 dido
X42 VDD VSS PCHG WREN SEL42 BL42 BL_42 DW42 DW_42 DR42 DR_42 dido
X43 VDD VSS PCHG WREN SEL43 BL43 BL_43 DW43 DW_43 DR43 DR_43 dido
X44 VDD VSS PCHG WREN SEL44 BL44 BL_44 DW44 DW_44 DR44 DR_44 dido
X45 VDD VSS PCHG WREN SEL45 BL45 BL_45 DW45 DW_45 DR45 DR_45 dido
X46 VDD VSS PCHG WREN SEL46 BL46 BL_46 DW46 DW_46 DR46 DR_46 dido
X47 VDD VSS PCHG WREN SEL47 BL47 BL_47 DW47 DW_47 DR47 DR_47 dido
X48 VDD VSS PCHG WREN SEL48 BL48 BL_48 DW48 DW_48 DR48 DR_48 dido
X49 VDD VSS PCHG WREN SEL49 BL49 BL_49 DW49 DW_49 DR49 DR_49 dido
X50 VDD VSS PCHG WREN SEL50 BL50 BL_50 DW50 DW_50 DR50 DR_50 dido
X51 VDD VSS PCHG WREN SEL51 BL51 BL_51 DW51 DW_51 DR51 DR_51 dido
X52 VDD VSS PCHG WREN SEL52 BL52 BL_52 DW52 DW_52 DR52 DR_52 dido
X53 VDD VSS PCHG WREN SEL53 BL53 BL_53 DW53 DW_53 DR53 DR_53 dido
X54 VDD VSS PCHG WREN SEL54 BL54 BL_54 DW54 DW_54 DR54 DR_54 dido
X55 VDD VSS PCHG WREN SEL55 BL55 BL_55 DW55 DW_55 DR55 DR_55 dido
X56 VDD VSS PCHG WREN SEL56 BL56 BL_56 DW56 DW_56 DR56 DR_56 dido
X57 VDD VSS PCHG WREN SEL57 BL57 BL_57 DW57 DW_57 DR57 DR_57 dido
X58 VDD VSS PCHG WREN SEL58 BL58 BL_58 DW58 DW_58 DR58 DR_58 dido
X59 VDD VSS PCHG WREN SEL59 BL59 BL_59 DW59 DW_59 DR59 DR_59 dido
X60 VDD VSS PCHG WREN SEL60 BL60 BL_60 DW60 DW_60 DR60 DR_60 dido
X61 VDD VSS PCHG WREN SEL61 BL61 BL_61 DW61 DW_61 DR61 DR_61 dido
X62 VDD VSS PCHG WREN SEL62 BL62 BL_62 DW62 DW_62 DR62 DR_62 dido
X63 VDD VSS PCHG WREN SEL63 BL63 BL_63 DW63 DW_63 DR63 DR_63 dido
.ends dido_arr_64

.subckt write_driver VDD VSS WREN Din DW DW_
X0 en_ WREN VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 en_ WREN VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X4 d_ Din VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X5 d_ Din VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X6 net1 Din VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X7 DW_ en_ net1 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X8 DW_ WREN net2 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
X9 net2 Din VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
X10 net3 d_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X11 DW en_ net3 VDD sky130_fd_pr__pfet_01v8 l=0.15 w=2
X12 DW WREN net4 VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
X13 net4 d_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=1
.ends write_driver

.subckt del10 VDD VSS A B
X0 VDD VSS A net1 notdel
X1 VDD VSS net1 net2 notdel
X2 VDD VSS net2 net3 notdel
X3 VDD VSS net3 net4 notdel
X4 VDD VSS net4 net5 notdel
X5 VDD VSS net5 net6 notdel
X6 VDD VSS net6 net7 notdel
X7 VDD VSS net7 net8 notdel
X8 VDD VSS net8 net9 notdel
X9 VDD VSS net9 net10 notdel
X10 VDD VSS net10 net11 notdel
X11 VDD VSS A net11 net12 nand2
X12 VDD VSS net12 B not
.ends del10

.subckt ctrl VDD VSS clk cs write DBL DBL_ WREN PCHG WLEN SAEN
X0 clk_ clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X1 clk_ clk VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X2 WLENP clk_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X3 WLENP clk_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=0.42
X4 VDD VSS write WREN_ not
X8 PCHG clk_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X9 PCHG clk_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
X10 DBL_ PCHG VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X11 DBL PCHG DBL_ VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X12 DBL PCHG VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=0.42
X13 VDD VSS cs WLENP WLENPP nand2
X21 WLEN WLENPP VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X22 WLEN WLENPP VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
X15 VDD VSS DBL_ RBL not
X16 VDD VSS WLEN RBL SAEN_ nand2
X17 SAEN SAEN_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X18 SAEN SAEN_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
X19 WREN WREN_ VDD VDD sky130_fd_pr__pfet_01v8 l=0.15 w=8
X20 WREN WREN_ VSS VSS sky130_fd_pr__nfet_01v8 l=0.15 w=4
.ends ctrl

.subckt input_reg8 VDD VSS clk D0 D1 D2 D3 D4 D5 D6 D7 Q0 Q1 Q2 Q3 Q4 Q5 Q6 Q7
X0 VDD VSS clk D0 Q0 in_reg
X1 VDD VSS clk D1 Q1 in_reg
X2 VDD VSS clk D2 Q2 in_reg
X3 VDD VSS clk D3 Q3 in_reg
X4 VDD VSS clk D4 Q4 in_reg
X5 VDD VSS clk D5 Q5 in_reg
X6 VDD VSS clk D6 Q6 in_reg
X7 VDD VSS clk D7 Q7 in_reg
.ends input_reg8

.subckt datain_reg64 VDD VSS clk WREN din0 din1 din2 din3 din4 din5 din6 din7 din8 din9 din10 din11 din12 din13 din14 din15 din16 din17 din18 din19 din20 din21 din22 din23 din24 din25 din26 din27 din28 din29 din30 din31 din32 din33 din34 din35 din36 din37 din38 din39 din40 din41 din42 din43 din44 din45 din46 din47 din48 din49 din50 din51 din52 din53 din54 din55 din56 din57 din58 din59 din60 din61 din62 din63 DW0 DW_0 DW1 DW_1 DW2 DW_2 DW3 DW_3 DW4 DW_4 DW5 DW_5 DW6 DW_6 DW7 DW_7 DW8 DW_8 DW9 DW_9 DW10 DW_10 DW11 DW_11 DW12 DW_12 DW13 DW_13 DW14 DW_14 DW15 DW_15 DW16 DW_16 DW17 DW_17 DW18 DW_18 DW19 DW_19 DW20 DW_20 DW21 DW_21 DW22 DW_22 DW23 DW_23 DW24 DW_24 DW25 DW_25 DW26 DW_26 DW27 DW_27 DW28 DW_28 DW29 DW_29 DW30 DW_30 DW31 DW_31 DW32 DW_32 DW33 DW_33 DW34 DW_34 DW35 DW_35 DW36 DW_36 DW37 DW_37 DW38 DW_38 DW39 DW_39 DW40 DW_40 DW41 DW_41 DW42 DW_42 DW43 DW_43 DW44 DW_44 DW45 DW_45 DW46 DW_46 DW47 DW_47 DW48 DW_48 DW49 DW_49 DW50 DW_50 DW51 DW_51 DW52 DW_52 DW53 DW_53 DW54 DW_54 DW55 DW_55 DW56 DW_56 DW57 DW_57 DW58 DW_58 DW59 DW_59 DW60 DW_60 DW61 DW_61 DW62 DW_62 DW63 DW_63
X0 VDD VSS clk din0 din_r0 in_reg
X1 VDD VSS clk din1 din_r1 in_reg
X2 VDD VSS clk din2 din_r2 in_reg
X3 VDD VSS clk din3 din_r3 in_reg
X4 VDD VSS clk din4 din_r4 in_reg
X5 VDD VSS clk din5 din_r5 in_reg
X6 VDD VSS clk din6 din_r6 in_reg
X7 VDD VSS clk din7 din_r7 in_reg
X8 VDD VSS clk din8 din_r8 in_reg
X9 VDD VSS clk din9 din_r9 in_reg
X10 VDD VSS clk din10 din_r10 in_reg
X11 VDD VSS clk din11 din_r11 in_reg
X12 VDD VSS clk din12 din_r12 in_reg
X13 VDD VSS clk din13 din_r13 in_reg
X14 VDD VSS clk din14 din_r14 in_reg
X15 VDD VSS clk din15 din_r15 in_reg
X16 VDD VSS clk din16 din_r16 in_reg
X17 VDD VSS clk din17 din_r17 in_reg
X18 VDD VSS clk din18 din_r18 in_reg
X19 VDD VSS clk din19 din_r19 in_reg
X20 VDD VSS clk din20 din_r20 in_reg
X21 VDD VSS clk din21 din_r21 in_reg
X22 VDD VSS clk din22 din_r22 in_reg
X23 VDD VSS clk din23 din_r23 in_reg
X24 VDD VSS clk din24 din_r24 in_reg
X25 VDD VSS clk din25 din_r25 in_reg
X26 VDD VSS clk din26 din_r26 in_reg
X27 VDD VSS clk din27 din_r27 in_reg
X28 VDD VSS clk din28 din_r28 in_reg
X29 VDD VSS clk din29 din_r29 in_reg
X30 VDD VSS clk din30 din_r30 in_reg
X31 VDD VSS clk din31 din_r31 in_reg
X32 VDD VSS clk din32 din_r32 in_reg
X33 VDD VSS clk din33 din_r33 in_reg
X34 VDD VSS clk din34 din_r34 in_reg
X35 VDD VSS clk din35 din_r35 in_reg
X36 VDD VSS clk din36 din_r36 in_reg
X37 VDD VSS clk din37 din_r37 in_reg
X38 VDD VSS clk din38 din_r38 in_reg
X39 VDD VSS clk din39 din_r39 in_reg
X40 VDD VSS clk din40 din_r40 in_reg
X41 VDD VSS clk din41 din_r41 in_reg
X42 VDD VSS clk din42 din_r42 in_reg
X43 VDD VSS clk din43 din_r43 in_reg
X44 VDD VSS clk din44 din_r44 in_reg
X45 VDD VSS clk din45 din_r45 in_reg
X46 VDD VSS clk din46 din_r46 in_reg
X47 VDD VSS clk din47 din_r47 in_reg
X48 VDD VSS clk din48 din_r48 in_reg
X49 VDD VSS clk din49 din_r49 in_reg
X50 VDD VSS clk din50 din_r50 in_reg
X51 VDD VSS clk din51 din_r51 in_reg
X52 VDD VSS clk din52 din_r52 in_reg
X53 VDD VSS clk din53 din_r53 in_reg
X54 VDD VSS clk din54 din_r54 in_reg
X55 VDD VSS clk din55 din_r55 in_reg
X56 VDD VSS clk din56 din_r56 in_reg
X57 VDD VSS clk din57 din_r57 in_reg
X58 VDD VSS clk din58 din_r58 in_reg
X59 VDD VSS clk din59 din_r59 in_reg
X60 VDD VSS clk din60 din_r60 in_reg
X61 VDD VSS clk din61 din_r61 in_reg
X62 VDD VSS clk din62 din_r62 in_reg
X63 VDD VSS clk din63 din_r63 in_reg
X64 VDD VSS WREN din_r0 DW0 DW_0 write_driver
X68 VDD VSS WREN din_r1 DW1 DW_1 write_driver
X72 VDD VSS WREN din_r2 DW2 DW_2 write_driver
X76 VDD VSS WREN din_r3 DW3 DW_3 write_driver
X80 VDD VSS WREN din_r4 DW4 DW_4 write_driver
X84 VDD VSS WREN din_r5 DW5 DW_5 write_driver
X88 VDD VSS WREN din_r6 DW6 DW_6 write_driver
X92 VDD VSS WREN din_r7 DW7 DW_7 write_driver
X96 VDD VSS WREN din_r8 DW8 DW_8 write_driver
X100 VDD VSS WREN din_r9 DW9 DW_9 write_driver
X104 VDD VSS WREN din_r10 DW10 DW_10 write_driver
X108 VDD VSS WREN din_r11 DW11 DW_11 write_driver
X112 VDD VSS WREN din_r12 DW12 DW_12 write_driver
X116 VDD VSS WREN din_r13 DW13 DW_13 write_driver
X120 VDD VSS WREN din_r14 DW14 DW_14 write_driver
X124 VDD VSS WREN din_r15 DW15 DW_15 write_driver
X128 VDD VSS WREN din_r16 DW16 DW_16 write_driver
X132 VDD VSS WREN din_r17 DW17 DW_17 write_driver
X136 VDD VSS WREN din_r18 DW18 DW_18 write_driver
X140 VDD VSS WREN din_r19 DW19 DW_19 write_driver
X144 VDD VSS WREN din_r20 DW20 DW_20 write_driver
X148 VDD VSS WREN din_r21 DW21 DW_21 write_driver
X152 VDD VSS WREN din_r22 DW22 DW_22 write_driver
X156 VDD VSS WREN din_r23 DW23 DW_23 write_driver
X160 VDD VSS WREN din_r24 DW24 DW_24 write_driver
X164 VDD VSS WREN din_r25 DW25 DW_25 write_driver
X168 VDD VSS WREN din_r26 DW26 DW_26 write_driver
X172 VDD VSS WREN din_r27 DW27 DW_27 write_driver
X176 VDD VSS WREN din_r28 DW28 DW_28 write_driver
X180 VDD VSS WREN din_r29 DW29 DW_29 write_driver
X184 VDD VSS WREN din_r30 DW30 DW_30 write_driver
X188 VDD VSS WREN din_r31 DW31 DW_31 write_driver
X192 VDD VSS WREN din_r32 DW32 DW_32 write_driver
X196 VDD VSS WREN din_r33 DW33 DW_33 write_driver
X200 VDD VSS WREN din_r34 DW34 DW_34 write_driver
X204 VDD VSS WREN din_r35 DW35 DW_35 write_driver
X208 VDD VSS WREN din_r36 DW36 DW_36 write_driver
X212 VDD VSS WREN din_r37 DW37 DW_37 write_driver
X216 VDD VSS WREN din_r38 DW38 DW_38 write_driver
X220 VDD VSS WREN din_r39 DW39 DW_39 write_driver
X224 VDD VSS WREN din_r40 DW40 DW_40 write_driver
X228 VDD VSS WREN din_r41 DW41 DW_41 write_driver
X232 VDD VSS WREN din_r42 DW42 DW_42 write_driver
X236 VDD VSS WREN din_r43 DW43 DW_43 write_driver
X240 VDD VSS WREN din_r44 DW44 DW_44 write_driver
X244 VDD VSS WREN din_r45 DW45 DW_45 write_driver
X248 VDD VSS WREN din_r46 DW46 DW_46 write_driver
X252 VDD VSS WREN din_r47 DW47 DW_47 write_driver
X256 VDD VSS WREN din_r48 DW48 DW_48 write_driver
X260 VDD VSS WREN din_r49 DW49 DW_49 write_driver
X264 VDD VSS WREN din_r50 DW50 DW_50 write_driver
X268 VDD VSS WREN din_r51 DW51 DW_51 write_driver
X272 VDD VSS WREN din_r52 DW52 DW_52 write_driver
X276 VDD VSS WREN din_r53 DW53 DW_53 write_driver
X280 VDD VSS WREN din_r54 DW54 DW_54 write_driver
X284 VDD VSS WREN din_r55 DW55 DW_55 write_driver
X288 VDD VSS WREN din_r56 DW56 DW_56 write_driver
X292 VDD VSS WREN din_r57 DW57 DW_57 write_driver
X296 VDD VSS WREN din_r58 DW58 DW_58 write_driver
X300 VDD VSS WREN din_r59 DW59 DW_59 write_driver
X304 VDD VSS WREN din_r60 DW60 DW_60 write_driver
X308 VDD VSS WREN din_r61 DW61 DW_61 write_driver
X312 VDD VSS WREN din_r62 DW62 DW_62 write_driver
X316 VDD VSS WREN din_r63 DW63 DW_63 write_driver
.ends datain_reg64

.subckt bit_arr_64 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL
X0 VDD VSS WL BL0 BL_0 bit_cell
X1 VDD VSS WL BL1 BL_1 bit_cell
X2 VDD VSS WL BL2 BL_2 bit_cell
X3 VDD VSS WL BL3 BL_3 bit_cell
X4 VDD VSS WL BL4 BL_4 bit_cell
X5 VDD VSS WL BL5 BL_5 bit_cell
X6 VDD VSS WL BL6 BL_6 bit_cell
X7 VDD VSS WL BL7 BL_7 bit_cell
X8 VDD VSS WL BL8 BL_8 bit_cell
X9 VDD VSS WL BL9 BL_9 bit_cell
X10 VDD VSS WL BL10 BL_10 bit_cell
X11 VDD VSS WL BL11 BL_11 bit_cell
X12 VDD VSS WL BL12 BL_12 bit_cell
X13 VDD VSS WL BL13 BL_13 bit_cell
X14 VDD VSS WL BL14 BL_14 bit_cell
X15 VDD VSS WL BL15 BL_15 bit_cell
X16 VDD VSS WL BL16 BL_16 bit_cell
X17 VDD VSS WL BL17 BL_17 bit_cell
X18 VDD VSS WL BL18 BL_18 bit_cell
X19 VDD VSS WL BL19 BL_19 bit_cell
X20 VDD VSS WL BL20 BL_20 bit_cell
X21 VDD VSS WL BL21 BL_21 bit_cell
X22 VDD VSS WL BL22 BL_22 bit_cell
X23 VDD VSS WL BL23 BL_23 bit_cell
X24 VDD VSS WL BL24 BL_24 bit_cell
X25 VDD VSS WL BL25 BL_25 bit_cell
X26 VDD VSS WL BL26 BL_26 bit_cell
X27 VDD VSS WL BL27 BL_27 bit_cell
X28 VDD VSS WL BL28 BL_28 bit_cell
X29 VDD VSS WL BL29 BL_29 bit_cell
X30 VDD VSS WL BL30 BL_30 bit_cell
X31 VDD VSS WL BL31 BL_31 bit_cell
X32 VDD VSS WL BL32 BL_32 bit_cell
X33 VDD VSS WL BL33 BL_33 bit_cell
X34 VDD VSS WL BL34 BL_34 bit_cell
X35 VDD VSS WL BL35 BL_35 bit_cell
X36 VDD VSS WL BL36 BL_36 bit_cell
X37 VDD VSS WL BL37 BL_37 bit_cell
X38 VDD VSS WL BL38 BL_38 bit_cell
X39 VDD VSS WL BL39 BL_39 bit_cell
X40 VDD VSS WL BL40 BL_40 bit_cell
X41 VDD VSS WL BL41 BL_41 bit_cell
X42 VDD VSS WL BL42 BL_42 bit_cell
X43 VDD VSS WL BL43 BL_43 bit_cell
X44 VDD VSS WL BL44 BL_44 bit_cell
X45 VDD VSS WL BL45 BL_45 bit_cell
X46 VDD VSS WL BL46 BL_46 bit_cell
X47 VDD VSS WL BL47 BL_47 bit_cell
X48 VDD VSS WL BL48 BL_48 bit_cell
X49 VDD VSS WL BL49 BL_49 bit_cell
X50 VDD VSS WL BL50 BL_50 bit_cell
X51 VDD VSS WL BL51 BL_51 bit_cell
X52 VDD VSS WL BL52 BL_52 bit_cell
X53 VDD VSS WL BL53 BL_53 bit_cell
X54 VDD VSS WL BL54 BL_54 bit_cell
X55 VDD VSS WL BL55 BL_55 bit_cell
X56 VDD VSS WL BL56 BL_56 bit_cell
X57 VDD VSS WL BL57 BL_57 bit_cell
X58 VDD VSS WL BL58 BL_58 bit_cell
X59 VDD VSS WL BL59 BL_59 bit_cell
X60 VDD VSS WL BL60 BL_60 bit_cell
X61 VDD VSS WL BL61 BL_61 bit_cell
X62 VDD VSS WL BL62 BL_62 bit_cell
X63 VDD VSS WL BL63 BL_63 bit_cell
.ends bit_arr_64

.subckt dmy_arr_128 VDD VSS WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 WL32 WL33 WL34 WL35 WL36 WL37 WL38 WL39 WL40 WL41 WL42 WL43 WL44 WL45 WL46 WL47 WL48 WL49 WL50 WL51 WL52 WL53 WL54 WL55 WL56 WL57 WL58 WL59 WL60 WL61 WL62 WL63 WL64 WL65 WL66 WL67 WL68 WL69 WL70 WL71 WL72 WL73 WL74 WL75 WL76 WL77 WL78 WL79 WL80 WL81 WL82 WL83 WL84 WL85 WL86 WL87 WL88 WL89 WL90 WL91 WL92 WL93 WL94 WL95 WL96 WL97 WL98 WL99 WL100 WL101 WL102 WL103 WL104 WL105 WL106 WL107 WL108 WL109 WL110 WL111 WL112 WL113 WL114 WL115 WL116 WL117 WL118 WL119 WL120 WL121 WL122 WL123 WL124 WL125 WL126 WL127 DBL DBL_
X0 VDD VSS WL0 DBL DBL_ dmy_cell
X1 VDD VSS WL1 DBL DBL_ dmy_cell
X2 VDD VSS WL2 DBL DBL_ dmy_cell
X3 VDD VSS WL3 DBL DBL_ dmy_cell
X4 VDD VSS WL4 DBL DBL_ dmy_cell
X5 VDD VSS WL5 DBL DBL_ dmy_cell
X6 VDD VSS WL6 DBL DBL_ dmy_cell
X7 VDD VSS WL7 DBL DBL_ dmy_cell
X8 VDD VSS WL8 DBL DBL_ dmy_cell
X9 VDD VSS WL9 DBL DBL_ dmy_cell
X10 VDD VSS WL10 DBL DBL_ dmy_cell
X11 VDD VSS WL11 DBL DBL_ dmy_cell
X12 VDD VSS WL12 DBL DBL_ dmy_cell
X13 VDD VSS WL13 DBL DBL_ dmy_cell
X14 VDD VSS WL14 DBL DBL_ dmy_cell
X15 VDD VSS WL15 DBL DBL_ dmy_cell
X16 VDD VSS WL16 DBL DBL_ dmy_cell
X17 VDD VSS WL17 DBL DBL_ dmy_cell
X18 VDD VSS WL18 DBL DBL_ dmy_cell
X19 VDD VSS WL19 DBL DBL_ dmy_cell
X20 VDD VSS WL20 DBL DBL_ dmy_cell
X21 VDD VSS WL21 DBL DBL_ dmy_cell
X22 VDD VSS WL22 DBL DBL_ dmy_cell
X23 VDD VSS WL23 DBL DBL_ dmy_cell
X24 VDD VSS WL24 DBL DBL_ dmy_cell
X25 VDD VSS WL25 DBL DBL_ dmy_cell
X26 VDD VSS WL26 DBL DBL_ dmy_cell
X27 VDD VSS WL27 DBL DBL_ dmy_cell
X28 VDD VSS WL28 DBL DBL_ dmy_cell
X29 VDD VSS WL29 DBL DBL_ dmy_cell
X30 VDD VSS WL30 DBL DBL_ dmy_cell
X31 VDD VSS WL31 DBL DBL_ dmy_cell
X32 VDD VSS WL32 DBL DBL_ dmy_cell
X33 VDD VSS WL33 DBL DBL_ dmy_cell
X34 VDD VSS WL34 DBL DBL_ dmy_cell
X35 VDD VSS WL35 DBL DBL_ dmy_cell
X36 VDD VSS WL36 DBL DBL_ dmy_cell
X37 VDD VSS WL37 DBL DBL_ dmy_cell
X38 VDD VSS WL38 DBL DBL_ dmy_cell
X39 VDD VSS WL39 DBL DBL_ dmy_cell
X40 VDD VSS WL40 DBL DBL_ dmy_cell
X41 VDD VSS WL41 DBL DBL_ dmy_cell
X42 VDD VSS WL42 DBL DBL_ dmy_cell
X43 VDD VSS WL43 DBL DBL_ dmy_cell
X44 VDD VSS WL44 DBL DBL_ dmy_cell
X45 VDD VSS WL45 DBL DBL_ dmy_cell
X46 VDD VSS WL46 DBL DBL_ dmy_cell
X47 VDD VSS WL47 DBL DBL_ dmy_cell
X48 VDD VSS WL48 DBL DBL_ dmy_cell
X49 VDD VSS WL49 DBL DBL_ dmy_cell
X50 VDD VSS WL50 DBL DBL_ dmy_cell
X51 VDD VSS WL51 DBL DBL_ dmy_cell
X52 VDD VSS WL52 DBL DBL_ dmy_cell
X53 VDD VSS WL53 DBL DBL_ dmy_cell
X54 VDD VSS WL54 DBL DBL_ dmy_cell
X55 VDD VSS WL55 DBL DBL_ dmy_cell
X56 VDD VSS WL56 DBL DBL_ dmy_cell
X57 VDD VSS WL57 DBL DBL_ dmy_cell
X58 VDD VSS WL58 DBL DBL_ dmy_cell
X59 VDD VSS WL59 DBL DBL_ dmy_cell
X60 VDD VSS WL60 DBL DBL_ dmy_cell
X61 VDD VSS WL61 DBL DBL_ dmy_cell
X62 VDD VSS WL62 DBL DBL_ dmy_cell
X63 VDD VSS WL63 DBL DBL_ dmy_cell
X64 VDD VSS WL64 DBL DBL_ dmy_cell
X65 VDD VSS WL65 DBL DBL_ dmy_cell
X66 VDD VSS WL66 DBL DBL_ dmy_cell
X67 VDD VSS WL67 DBL DBL_ dmy_cell
X68 VDD VSS WL68 DBL DBL_ dmy_cell
X69 VDD VSS WL69 DBL DBL_ dmy_cell
X70 VDD VSS WL70 DBL DBL_ dmy_cell
X71 VDD VSS WL71 DBL DBL_ dmy_cell
X72 VDD VSS WL72 DBL DBL_ dmy_cell
X73 VDD VSS WL73 DBL DBL_ dmy_cell
X74 VDD VSS WL74 DBL DBL_ dmy_cell
X75 VDD VSS WL75 DBL DBL_ dmy_cell
X76 VDD VSS WL76 DBL DBL_ dmy_cell
X77 VDD VSS WL77 DBL DBL_ dmy_cell
X78 VDD VSS WL78 DBL DBL_ dmy_cell
X79 VDD VSS WL79 DBL DBL_ dmy_cell
X80 VDD VSS WL80 DBL DBL_ dmy_cell
X81 VDD VSS WL81 DBL DBL_ dmy_cell
X82 VDD VSS WL82 DBL DBL_ dmy_cell
X83 VDD VSS WL83 DBL DBL_ dmy_cell
X84 VDD VSS WL84 DBL DBL_ dmy_cell
X85 VDD VSS WL85 DBL DBL_ dmy_cell
X86 VDD VSS WL86 DBL DBL_ dmy_cell
X87 VDD VSS WL87 DBL DBL_ dmy_cell
X88 VDD VSS WL88 DBL DBL_ dmy_cell
X89 VDD VSS WL89 DBL DBL_ dmy_cell
X90 VDD VSS WL90 DBL DBL_ dmy_cell
X91 VDD VSS WL91 DBL DBL_ dmy_cell
X92 VDD VSS WL92 DBL DBL_ dmy_cell
X93 VDD VSS WL93 DBL DBL_ dmy_cell
X94 VDD VSS WL94 DBL DBL_ dmy_cell
X95 VDD VSS WL95 DBL DBL_ dmy_cell
X96 VDD VSS WL96 DBL DBL_ dmy_cell
X97 VDD VSS WL97 DBL DBL_ dmy_cell
X98 VDD VSS WL98 DBL DBL_ dmy_cell
X99 VDD VSS WL99 DBL DBL_ dmy_cell
X100 VDD VSS WL100 DBL DBL_ dmy_cell
X101 VDD VSS WL101 DBL DBL_ dmy_cell
X102 VDD VSS WL102 DBL DBL_ dmy_cell
X103 VDD VSS WL103 DBL DBL_ dmy_cell
X104 VDD VSS WL104 DBL DBL_ dmy_cell
X105 VDD VSS WL105 DBL DBL_ dmy_cell
X106 VDD VSS WL106 DBL DBL_ dmy_cell
X107 VDD VSS WL107 DBL DBL_ dmy_cell
X108 VDD VSS WL108 DBL DBL_ dmy_cell
X109 VDD VSS WL109 DBL DBL_ dmy_cell
X110 VDD VSS WL110 DBL DBL_ dmy_cell
X111 VDD VSS WL111 DBL DBL_ dmy_cell
X112 VDD VSS WL112 DBL DBL_ dmy_cell
X113 VDD VSS WL113 DBL DBL_ dmy_cell
X114 VDD VSS WL114 DBL DBL_ dmy_cell
X115 VDD VSS WL115 DBL DBL_ dmy_cell
X116 VDD VSS WL116 DBL DBL_ dmy_cell
X117 VDD VSS WL117 DBL DBL_ dmy_cell
X118 VDD VSS WL118 DBL DBL_ dmy_cell
X119 VDD VSS WL119 DBL DBL_ dmy_cell
X120 VDD VSS WL120 DBL DBL_ dmy_cell
X121 VDD VSS WL121 DBL DBL_ dmy_cell
X122 VDD VSS WL122 DBL DBL_ dmy_cell
X123 VDD VSS WL123 DBL DBL_ dmy_cell
X124 VDD VSS WL124 DBL DBL_ dmy_cell
X125 VDD VSS WL125 DBL DBL_ dmy_cell
X126 VDD VSS WL126 DBL DBL_ dmy_cell
X127 VDD VSS WL127 DBL DBL_ dmy_cell
.ends dmy_arr_128

.subckt se_arr_64 VDD VSS SAEN BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 SB0 SB1 SB2 SB3 SB4 SB5 SB6 SB7 SB8 SB9 SB10 SB11 SB12 SB13 SB14 SB15 SB16 SB17 SB18 SB19 SB20 SB21 SB22 SB23 SB24 SB25 SB26 SB27 SB28 SB29 SB30 SB31 SB32 SB33 SB34 SB35 SB36 SB37 SB38 SB39 SB40 SB41 SB42 SB43 SB44 SB45 SB46 SB47 SB48 SB49 SB50 SB51 SB52 SB53 SB54 SB55 SB56 SB57 SB58 SB59 SB60 SB61 SB62 SB63
X0 VDD VSS SAEN BL0 BL_0 SB0 se_cell
X1 VDD VSS SAEN BL1 BL_1 SB1 se_cell
X2 VDD VSS SAEN BL2 BL_2 SB2 se_cell
X3 VDD VSS SAEN BL3 BL_3 SB3 se_cell
X4 VDD VSS SAEN BL4 BL_4 SB4 se_cell
X5 VDD VSS SAEN BL5 BL_5 SB5 se_cell
X6 VDD VSS SAEN BL6 BL_6 SB6 se_cell
X7 VDD VSS SAEN BL7 BL_7 SB7 se_cell
X8 VDD VSS SAEN BL8 BL_8 SB8 se_cell
X9 VDD VSS SAEN BL9 BL_9 SB9 se_cell
X10 VDD VSS SAEN BL10 BL_10 SB10 se_cell
X11 VDD VSS SAEN BL11 BL_11 SB11 se_cell
X12 VDD VSS SAEN BL12 BL_12 SB12 se_cell
X13 VDD VSS SAEN BL13 BL_13 SB13 se_cell
X14 VDD VSS SAEN BL14 BL_14 SB14 se_cell
X15 VDD VSS SAEN BL15 BL_15 SB15 se_cell
X16 VDD VSS SAEN BL16 BL_16 SB16 se_cell
X17 VDD VSS SAEN BL17 BL_17 SB17 se_cell
X18 VDD VSS SAEN BL18 BL_18 SB18 se_cell
X19 VDD VSS SAEN BL19 BL_19 SB19 se_cell
X20 VDD VSS SAEN BL20 BL_20 SB20 se_cell
X21 VDD VSS SAEN BL21 BL_21 SB21 se_cell
X22 VDD VSS SAEN BL22 BL_22 SB22 se_cell
X23 VDD VSS SAEN BL23 BL_23 SB23 se_cell
X24 VDD VSS SAEN BL24 BL_24 SB24 se_cell
X25 VDD VSS SAEN BL25 BL_25 SB25 se_cell
X26 VDD VSS SAEN BL26 BL_26 SB26 se_cell
X27 VDD VSS SAEN BL27 BL_27 SB27 se_cell
X28 VDD VSS SAEN BL28 BL_28 SB28 se_cell
X29 VDD VSS SAEN BL29 BL_29 SB29 se_cell
X30 VDD VSS SAEN BL30 BL_30 SB30 se_cell
X31 VDD VSS SAEN BL31 BL_31 SB31 se_cell
X32 VDD VSS SAEN BL32 BL_32 SB32 se_cell
X33 VDD VSS SAEN BL33 BL_33 SB33 se_cell
X34 VDD VSS SAEN BL34 BL_34 SB34 se_cell
X35 VDD VSS SAEN BL35 BL_35 SB35 se_cell
X36 VDD VSS SAEN BL36 BL_36 SB36 se_cell
X37 VDD VSS SAEN BL37 BL_37 SB37 se_cell
X38 VDD VSS SAEN BL38 BL_38 SB38 se_cell
X39 VDD VSS SAEN BL39 BL_39 SB39 se_cell
X40 VDD VSS SAEN BL40 BL_40 SB40 se_cell
X41 VDD VSS SAEN BL41 BL_41 SB41 se_cell
X42 VDD VSS SAEN BL42 BL_42 SB42 se_cell
X43 VDD VSS SAEN BL43 BL_43 SB43 se_cell
X44 VDD VSS SAEN BL44 BL_44 SB44 se_cell
X45 VDD VSS SAEN BL45 BL_45 SB45 se_cell
X46 VDD VSS SAEN BL46 BL_46 SB46 se_cell
X47 VDD VSS SAEN BL47 BL_47 SB47 se_cell
X48 VDD VSS SAEN BL48 BL_48 SB48 se_cell
X49 VDD VSS SAEN BL49 BL_49 SB49 se_cell
X50 VDD VSS SAEN BL50 BL_50 SB50 se_cell
X51 VDD VSS SAEN BL51 BL_51 SB51 se_cell
X52 VDD VSS SAEN BL52 BL_52 SB52 se_cell
X53 VDD VSS SAEN BL53 BL_53 SB53 se_cell
X54 VDD VSS SAEN BL54 BL_54 SB54 se_cell
X55 VDD VSS SAEN BL55 BL_55 SB55 se_cell
X56 VDD VSS SAEN BL56 BL_56 SB56 se_cell
X57 VDD VSS SAEN BL57 BL_57 SB57 se_cell
X58 VDD VSS SAEN BL58 BL_58 SB58 se_cell
X59 VDD VSS SAEN BL59 BL_59 SB59 se_cell
X60 VDD VSS SAEN BL60 BL_60 SB60 se_cell
X61 VDD VSS SAEN BL61 BL_61 SB61 se_cell
X62 VDD VSS SAEN BL62 BL_62 SB62 se_cell
X63 VDD VSS SAEN BL63 BL_63 SB63 se_cell
.ends se_arr_64

.subckt mat_arr_64 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 WL32 WL33 WL34 WL35 WL36 WL37 WL38 WL39 WL40 WL41 WL42 WL43 WL44 WL45 WL46 WL47 WL48 WL49 WL50 WL51 WL52 WL53 WL54 WL55 WL56 WL57 WL58 WL59 WL60 WL61 WL62 WL63 WL64 WL65 WL66 WL67 WL68 WL69 WL70 WL71 WL72 WL73 WL74 WL75 WL76 WL77 WL78 WL79 WL80 WL81 WL82 WL83 WL84 WL85 WL86 WL87 WL88 WL89 WL90 WL91 WL92 WL93 WL94 WL95 WL96 WL97 WL98 WL99 WL100 WL101 WL102 WL103 WL104 WL105 WL106 WL107 WL108 WL109 WL110 WL111 WL112 WL113 WL114 WL115 WL116 WL117 WL118 WL119 WL120 WL121 WL122 WL123 WL124 WL125 WL126 WL127
X0 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL0 bit_arr_64
X1 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL1 bit_arr_64
X2 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL2 bit_arr_64
X3 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL3 bit_arr_64
X4 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL4 bit_arr_64
X5 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL5 bit_arr_64
X6 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL6 bit_arr_64
X7 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL7 bit_arr_64
X8 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL8 bit_arr_64
X9 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL9 bit_arr_64
X10 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL10 bit_arr_64
X11 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL11 bit_arr_64
X12 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL12 bit_arr_64
X13 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL13 bit_arr_64
X14 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL14 bit_arr_64
X15 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL15 bit_arr_64
X16 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL16 bit_arr_64
X17 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL17 bit_arr_64
X18 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL18 bit_arr_64
X19 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL19 bit_arr_64
X20 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL20 bit_arr_64
X21 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL21 bit_arr_64
X22 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL22 bit_arr_64
X23 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL23 bit_arr_64
X24 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL24 bit_arr_64
X25 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL25 bit_arr_64
X26 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL26 bit_arr_64
X27 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL27 bit_arr_64
X28 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL28 bit_arr_64
X29 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL29 bit_arr_64
X30 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL30 bit_arr_64
X31 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL31 bit_arr_64
X32 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL32 bit_arr_64
X33 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL33 bit_arr_64
X34 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL34 bit_arr_64
X35 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL35 bit_arr_64
X36 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL36 bit_arr_64
X37 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL37 bit_arr_64
X38 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL38 bit_arr_64
X39 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL39 bit_arr_64
X40 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL40 bit_arr_64
X41 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL41 bit_arr_64
X42 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL42 bit_arr_64
X43 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL43 bit_arr_64
X44 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL44 bit_arr_64
X45 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL45 bit_arr_64
X46 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL46 bit_arr_64
X47 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL47 bit_arr_64
X48 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL48 bit_arr_64
X49 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL49 bit_arr_64
X50 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL50 bit_arr_64
X51 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL51 bit_arr_64
X52 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL52 bit_arr_64
X53 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL53 bit_arr_64
X54 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL54 bit_arr_64
X55 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL55 bit_arr_64
X56 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL56 bit_arr_64
X57 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL57 bit_arr_64
X58 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL58 bit_arr_64
X59 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL59 bit_arr_64
X60 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL60 bit_arr_64
X61 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL61 bit_arr_64
X62 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL62 bit_arr_64
X63 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL63 bit_arr_64
X64 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL64 bit_arr_64
X65 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL65 bit_arr_64
X66 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL66 bit_arr_64
X67 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL67 bit_arr_64
X68 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL68 bit_arr_64
X69 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL69 bit_arr_64
X70 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL70 bit_arr_64
X71 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL71 bit_arr_64
X72 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL72 bit_arr_64
X73 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL73 bit_arr_64
X74 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL74 bit_arr_64
X75 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL75 bit_arr_64
X76 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL76 bit_arr_64
X77 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL77 bit_arr_64
X78 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL78 bit_arr_64
X79 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL79 bit_arr_64
X80 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL80 bit_arr_64
X81 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL81 bit_arr_64
X82 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL82 bit_arr_64
X83 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL83 bit_arr_64
X84 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL84 bit_arr_64
X85 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL85 bit_arr_64
X86 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL86 bit_arr_64
X87 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL87 bit_arr_64
X88 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL88 bit_arr_64
X89 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL89 bit_arr_64
X90 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL90 bit_arr_64
X91 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL91 bit_arr_64
X92 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL92 bit_arr_64
X93 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL93 bit_arr_64
X94 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL94 bit_arr_64
X95 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL95 bit_arr_64
X96 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL96 bit_arr_64
X97 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL97 bit_arr_64
X98 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL98 bit_arr_64
X99 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL99 bit_arr_64
X100 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL100 bit_arr_64
X101 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL101 bit_arr_64
X102 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL102 bit_arr_64
X103 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL103 bit_arr_64
X104 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL104 bit_arr_64
X105 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL105 bit_arr_64
X106 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL106 bit_arr_64
X107 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL107 bit_arr_64
X108 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL108 bit_arr_64
X109 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL109 bit_arr_64
X110 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL110 bit_arr_64
X111 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL111 bit_arr_64
X112 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL112 bit_arr_64
X113 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL113 bit_arr_64
X114 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL114 bit_arr_64
X115 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL115 bit_arr_64
X116 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL116 bit_arr_64
X117 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL117 bit_arr_64
X118 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL118 bit_arr_64
X119 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL119 bit_arr_64
X120 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL120 bit_arr_64
X121 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL121 bit_arr_64
X122 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL122 bit_arr_64
X123 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL123 bit_arr_64
X124 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL124 bit_arr_64
X125 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL125 bit_arr_64
X126 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL126 bit_arr_64
X127 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL127 bit_arr_64
.ends mat_arr_64

.subckt sram128x64 VDD VSS clk addr0 addr1 addr2 addr3 addr4 addr5 addr6 din0 din1 din2 din3 din4 din5 din6 din7 din8 din9 din10 din11 din12 din13 din14 din15 din16 din17 din18 din19 din20 din21 din22 din23 din24 din25 din26 din27 din28 din29 din30 din31 din32 din33 din34 din35 din36 din37 din38 din39 din40 din41 din42 din43 din44 din45 din46 din47 din48 din49 din50 din51 din52 din53 din54 din55 din56 din57 din58 din59 din60 din61 din62 din63 Q0 Q1 Q2 Q3 Q4 Q5 Q6 Q7 Q8 Q9 Q10 Q11 Q12 Q13 Q14 Q15 Q16 Q17 Q18 Q19 Q20 Q21 Q22 Q23 Q24 Q25 Q26 Q27 Q28 Q29 Q30 Q31 Q32 Q33 Q34 Q35 Q36 Q37 Q38 Q39 Q40 Q41 Q42 Q43 Q44 Q45 Q46 Q47 Q48 Q49 Q50 Q51 Q52 Q53 Q54 Q55 Q56 Q57 Q58 Q59 Q60 Q61 Q62 Q63 w_en cs
X0 VDD VSS clk addr0 addr1 addr2 addr3 addr4 addr5 addr6 w_en A0 A1 A2 A3 A4 A5 A6 write input_reg8
X1 VDD VSS A0 A1 A2 A3 A4 A5 A6 DC0 DC1 DC2 DC3 DC4 DC5 DC6 DC7 DC8 DC9 DC10 DC11 DC12 DC13 DC14 DC15 DC16 DC17 DC18 DC19 DC20 DC21 DC22 DC23 DC24 DC25 DC26 DC27 DC28 DC29 DC30 DC31 DC32 DC33 DC34 DC35 DC36 DC37 DC38 DC39 DC40 DC41 DC42 DC43 DC44 DC45 DC46 DC47 DC48 DC49 DC50 DC51 DC52 DC53 DC54 DC55 DC56 DC57 DC58 DC59 DC60 DC61 DC62 DC63 DC64 DC65 DC66 DC67 DC68 DC69 DC70 DC71 DC72 DC73 DC74 DC75 DC76 DC77 DC78 DC79 DC80 DC81 DC82 DC83 DC84 DC85 DC86 DC87 DC88 DC89 DC90 DC91 DC92 DC93 DC94 DC95 DC96 DC97 DC98 DC99 DC100 DC101 DC102 DC103 DC104 DC105 DC106 DC107 DC108 DC109 DC110 DC111 DC112 DC113 DC114 DC115 DC116 DC117 DC118 DC119 DC120 DC121 DC122 DC123 DC124 DC125 DC126 DC127 row_dec128
X2 VDD VSS WLEN DC0 DC1 DC2 DC3 DC4 DC5 DC6 DC7 DC8 DC9 DC10 DC11 DC12 DC13 DC14 DC15 DC16 DC17 DC18 DC19 DC20 DC21 DC22 DC23 DC24 DC25 DC26 DC27 DC28 DC29 DC30 DC31 DC32 DC33 DC34 DC35 DC36 DC37 DC38 DC39 DC40 DC41 DC42 DC43 DC44 DC45 DC46 DC47 DC48 DC49 DC50 DC51 DC52 DC53 DC54 DC55 DC56 DC57 DC58 DC59 DC60 DC61 DC62 DC63 DC64 DC65 DC66 DC67 DC68 DC69 DC70 DC71 DC72 DC73 DC74 DC75 DC76 DC77 DC78 DC79 DC80 DC81 DC82 DC83 DC84 DC85 DC86 DC87 DC88 DC89 DC90 DC91 DC92 DC93 DC94 DC95 DC96 DC97 DC98 DC99 DC100 DC101 DC102 DC103 DC104 DC105 DC106 DC107 DC108 DC109 DC110 DC111 DC112 DC113 DC114 DC115 DC116 DC117 DC118 DC119 DC120 DC121 DC122 DC123 DC124 DC125 DC126 DC127 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 WL32 WL33 WL34 WL35 WL36 WL37 WL38 WL39 WL40 WL41 WL42 WL43 WL44 WL45 WL46 WL47 WL48 WL49 WL50 WL51 WL52 WL53 WL54 WL55 WL56 WL57 WL58 WL59 WL60 WL61 WL62 WL63 WL64 WL65 WL66 WL67 WL68 WL69 WL70 WL71 WL72 WL73 WL74 WL75 WL76 WL77 WL78 WL79 WL80 WL81 WL82 WL83 WL84 WL85 WL86 WL87 WL88 WL89 WL90 WL91 WL92 WL93 WL94 WL95 WL96 WL97 WL98 WL99 WL100 WL101 WL102 WL103 WL104 WL105 WL106 WL107 WL108 WL109 WL110 WL111 WL112 WL113 WL114 WL115 WL116 WL117 WL118 WL119 WL120 WL121 WL122 WL123 WL124 WL125 WL126 WL127 rd_arr_128
X3 VDD VSS WLEN SEL0 not
X4 VDD VSS PCHG WREN SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 SEL0 BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 DW0 DW_0 DW1 DW_1 DW2 DW_2 DW3 DW_3 DW4 DW_4 DW5 DW_5 DW6 DW_6 DW7 DW_7 DW8 DW_8 DW9 DW_9 DW10 DW_10 DW11 DW_11 DW12 DW_12 DW13 DW_13 DW14 DW_14 DW15 DW_15 DW16 DW_16 DW17 DW_17 DW18 DW_18 DW19 DW_19 DW20 DW_20 DW21 DW_21 DW22 DW_22 DW23 DW_23 DW24 DW_24 DW25 DW_25 DW26 DW_26 DW27 DW_27 DW28 DW_28 DW29 DW_29 DW30 DW_30 DW31 DW_31 DW32 DW_32 DW33 DW_33 DW34 DW_34 DW35 DW_35 DW36 DW_36 DW37 DW_37 DW38 DW_38 DW39 DW_39 DW40 DW_40 DW41 DW_41 DW42 DW_42 DW43 DW_43 DW44 DW_44 DW45 DW_45 DW46 DW_46 DW47 DW_47 DW48 DW_48 DW49 DW_49 DW50 DW_50 DW51 DW_51 DW52 DW_52 DW53 DW_53 DW54 DW_54 DW55 DW_55 DW56 DW_56 DW57 DW_57 DW58 DW_58 DW59 DW_59 DW60 DW_60 DW61 DW_61 DW62 DW_62 DW63 DW_63 DR0 DR_0 DR1 DR_1 DR2 DR_2 DR3 DR_3 DR4 DR_4 DR5 DR_5 DR6 DR_6 DR7 DR_7 DR8 DR_8 DR9 DR_9 DR10 DR_10 DR11 DR_11 DR12 DR_12 DR13 DR_13 DR14 DR_14 DR15 DR_15 DR16 DR_16 DR17 DR_17 DR18 DR_18 DR19 DR_19 DR20 DR_20 DR21 DR_21 DR22 DR_22 DR23 DR_23 DR24 DR_24 DR25 DR_25 DR26 DR_26 DR27 DR_27 DR28 DR_28 DR29 DR_29 DR30 DR_30 DR31 DR_31 DR32 DR_32 DR33 DR_33 DR34 DR_34 DR35 DR_35 DR36 DR_36 DR37 DR_37 DR38 DR_38 DR39 DR_39 DR40 DR_40 DR41 DR_41 DR42 DR_42 DR43 DR_43 DR44 DR_44 DR45 DR_45 DR46 DR_46 DR47 DR_47 DR48 DR_48 DR49 DR_49 DR50 DR_50 DR51 DR_51 DR52 DR_52 DR53 DR_53 DR54 DR_54 DR55 DR_55 DR56 DR_56 DR57 DR_57 DR58 DR_58 DR59 DR_59 DR60 DR_60 DR61 DR_61 DR62 DR_62 DR63 DR_63 dido_arr_64
X5 VDD VSS clk WREN din0 din1 din2 din3 din4 din5 din6 din7 din8 din9 din10 din11 din12 din13 din14 din15 din16 din17 din18 din19 din20 din21 din22 din23 din24 din25 din26 din27 din28 din29 din30 din31 din32 din33 din34 din35 din36 din37 din38 din39 din40 din41 din42 din43 din44 din45 din46 din47 din48 din49 din50 din51 din52 din53 din54 din55 din56 din57 din58 din59 din60 din61 din62 din63 DW0 DW_0 DW1 DW_1 DW2 DW_2 DW3 DW_3 DW4 DW_4 DW5 DW_5 DW6 DW_6 DW7 DW_7 DW8 DW_8 DW9 DW_9 DW10 DW_10 DW11 DW_11 DW12 DW_12 DW13 DW_13 DW14 DW_14 DW15 DW_15 DW16 DW_16 DW17 DW_17 DW18 DW_18 DW19 DW_19 DW20 DW_20 DW21 DW_21 DW22 DW_22 DW23 DW_23 DW24 DW_24 DW25 DW_25 DW26 DW_26 DW27 DW_27 DW28 DW_28 DW29 DW_29 DW30 DW_30 DW31 DW_31 DW32 DW_32 DW33 DW_33 DW34 DW_34 DW35 DW_35 DW36 DW_36 DW37 DW_37 DW38 DW_38 DW39 DW_39 DW40 DW_40 DW41 DW_41 DW42 DW_42 DW43 DW_43 DW44 DW_44 DW45 DW_45 DW46 DW_46 DW47 DW_47 DW48 DW_48 DW49 DW_49 DW50 DW_50 DW51 DW_51 DW52 DW_52 DW53 DW_53 DW54 DW_54 DW55 DW_55 DW56 DW_56 DW57 DW_57 DW58 DW_58 DW59 DW_59 DW60 DW_60 DW61 DW_61 DW62 DW_62 DW63 DW_63 datain_reg64
X6 VDD VSS BL0 BL_0 BL1 BL_1 BL2 BL_2 BL3 BL_3 BL4 BL_4 BL5 BL_5 BL6 BL_6 BL7 BL_7 BL8 BL_8 BL9 BL_9 BL10 BL_10 BL11 BL_11 BL12 BL_12 BL13 BL_13 BL14 BL_14 BL15 BL_15 BL16 BL_16 BL17 BL_17 BL18 BL_18 BL19 BL_19 BL20 BL_20 BL21 BL_21 BL22 BL_22 BL23 BL_23 BL24 BL_24 BL25 BL_25 BL26 BL_26 BL27 BL_27 BL28 BL_28 BL29 BL_29 BL30 BL_30 BL31 BL_31 BL32 BL_32 BL33 BL_33 BL34 BL_34 BL35 BL_35 BL36 BL_36 BL37 BL_37 BL38 BL_38 BL39 BL_39 BL40 BL_40 BL41 BL_41 BL42 BL_42 BL43 BL_43 BL44 BL_44 BL45 BL_45 BL46 BL_46 BL47 BL_47 BL48 BL_48 BL49 BL_49 BL50 BL_50 BL51 BL_51 BL52 BL_52 BL53 BL_53 BL54 BL_54 BL55 BL_55 BL56 BL_56 BL57 BL_57 BL58 BL_58 BL59 BL_59 BL60 BL_60 BL61 BL_61 BL62 BL_62 BL63 BL_63 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 WL32 WL33 WL34 WL35 WL36 WL37 WL38 WL39 WL40 WL41 WL42 WL43 WL44 WL45 WL46 WL47 WL48 WL49 WL50 WL51 WL52 WL53 WL54 WL55 WL56 WL57 WL58 WL59 WL60 WL61 WL62 WL63 WL64 WL65 WL66 WL67 WL68 WL69 WL70 WL71 WL72 WL73 WL74 WL75 WL76 WL77 WL78 WL79 WL80 WL81 WL82 WL83 WL84 WL85 WL86 WL87 WL88 WL89 WL90 WL91 WL92 WL93 WL94 WL95 WL96 WL97 WL98 WL99 WL100 WL101 WL102 WL103 WL104 WL105 WL106 WL107 WL108 WL109 WL110 WL111 WL112 WL113 WL114 WL115 WL116 WL117 WL118 WL119 WL120 WL121 WL122 WL123 WL124 WL125 WL126 WL127 mat_arr_64
X7 VDD VSS SAEN DR0 DR_0 DR1 DR_1 DR2 DR_2 DR3 DR_3 DR4 DR_4 DR5 DR_5 DR6 DR_6 DR7 DR_7 DR8 DR_8 DR9 DR_9 DR10 DR_10 DR11 DR_11 DR12 DR_12 DR13 DR_13 DR14 DR_14 DR15 DR_15 DR16 DR_16 DR17 DR_17 DR18 DR_18 DR19 DR_19 DR20 DR_20 DR21 DR_21 DR22 DR_22 DR23 DR_23 DR24 DR_24 DR25 DR_25 DR26 DR_26 DR27 DR_27 DR28 DR_28 DR29 DR_29 DR30 DR_30 DR31 DR_31 DR32 DR_32 DR33 DR_33 DR34 DR_34 DR35 DR_35 DR36 DR_36 DR37 DR_37 DR38 DR_38 DR39 DR_39 DR40 DR_40 DR41 DR_41 DR42 DR_42 DR43 DR_43 DR44 DR_44 DR45 DR_45 DR46 DR_46 DR47 DR_47 DR48 DR_48 DR49 DR_49 DR50 DR_50 DR51 DR_51 DR52 DR_52 DR53 DR_53 DR54 DR_54 DR55 DR_55 DR56 DR_56 DR57 DR_57 DR58 DR_58 DR59 DR_59 DR60 DR_60 DR61 DR_61 DR62 DR_62 DR63 DR_63 Q0 Q1 Q2 Q3 Q4 Q5 Q6 Q7 Q8 Q9 Q10 Q11 Q12 Q13 Q14 Q15 Q16 Q17 Q18 Q19 Q20 Q21 Q22 Q23 Q24 Q25 Q26 Q27 Q28 Q29 Q30 Q31 Q32 Q33 Q34 Q35 Q36 Q37 Q38 Q39 Q40 Q41 Q42 Q43 Q44 Q45 Q46 Q47 Q48 Q49 Q50 Q51 Q52 Q53 Q54 Q55 Q56 Q57 Q58 Q59 Q60 Q61 Q62 Q63 se_arr_64
X8 VDD VSS clk cs write DBL DBL_ WREN PCHG WLEN SAEN ctrl
X9 VDD VSS WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16 WL17 WL18 WL19 WL20 WL21 WL22 WL23 WL24 WL25 WL26 WL27 WL28 WL29 WL30 WL31 WL32 WL33 WL34 WL35 WL36 WL37 WL38 WL39 WL40 WL41 WL42 WL43 WL44 WL45 WL46 WL47 WL48 WL49 WL50 WL51 WL52 WL53 WL54 WL55 WL56 WL57 WL58 WL59 WL60 WL61 WL62 WL63 WL64 WL65 WL66 WL67 WL68 WL69 WL70 WL71 WL72 WL73 WL74 WL75 WL76 WL77 WL78 WL79 WL80 WL81 WL82 WL83 WL84 WL85 WL86 WL87 WL88 WL89 WL90 WL91 WL92 WL93 WL94 WL95 WL96 WL97 WL98 WL99 WL100 WL101 WL102 WL103 WL104 WL105 WL106 WL107 WL108 WL109 WL110 WL111 WL112 WL113 WL114 WL115 WL116 WL117 WL118 WL119 WL120 WL121 WL122 WL123 WL124 WL125 WL126 WL127 DBL DBL_ dmy_arr_128
.ends sram128x64

