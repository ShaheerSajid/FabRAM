.title characterizer
.include /home/shaheer/Desktop/FabRAM/FE/out/sram32x4.spi
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

      .tran 0.01194755n 23.8951n 11.94755n
      .control
      set hcopydevtype = svg
      run
      meas tran tdiff_cell_rise TRIG v(clk) VAL=0.9 RISE=1 TARG v(Q0) VAL=0.9 RISE=1 
      meas tran tdiff_tran_rise TRIG v(Q0)  VAL=0.18000000000000002 RISE=1 TARG v(Q0) VAL=1.62 RISE=1 
      meas tran tdiff_cell_fall TRIG v(clk) VAL=0.9 RISE=2 TARG v(Q0) VAL=0.9 FALL=1 
      meas tran tdiff_tran_fall TRIG v(Q0)  VAL=1.62 FALL=1 TARG v(Q0) VAL=0.18000000000000002 FALL=1 

      echo "$&tdiff_cell_rise,$&tdiff_tran_rise $&tdiff_cell_fall,$&tdiff_tran_fall" > log/sim_0.38951_0.03289.text
      hardcopy log/sim_0.38951_0.03289.svg v(clk) v(Q0) v(x0.PCHG) v(x0.WLEN) v(x0.SAEN) v(x0.x8.RSTP)
      exit
      .endc
      
Vpower VDD 0 1.8
Vgnd VSS 0 0
Vclk clk VSS DC 0V PULSE(0V 1.8V 0ns 0.48688750000000003ns 0.48688750000000003ns 2.5ns 5.973775ns)
Vaddr addr VSS DC 0V PULSE(0V 1.8V 0s 1ps 1ps 2.5ns 11.94755ns)
Vdin din VSS DC 0V PULSE(0V 1.8V 0s 1ps 1ps 2.5ns 11.94755ns)
Vwrite write VSS DC 0V PULSE(0V 1.8V 0s 1ps 1ps 11.94755ns 23.8951ns)
X0 VDD VSS clk addr addr addr addr addr din din din din Q0 Q1 Q2 Q3 write sram32x4
C0 Q0 VSS 0.03289p
