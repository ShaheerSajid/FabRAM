magic
tech sky130A
magscale 1 2
timestamp 1702464972
<< poly >>
rect 94 472 124 477
rect 44 456 124 472
rect 44 422 60 456
rect 94 422 124 456
rect 44 406 124 422
rect 94 264 124 406
rect 182 400 212 477
rect 170 384 224 400
rect 170 350 180 384
rect 214 350 224 384
rect 170 334 224 350
rect 182 263 212 334
rect 270 326 300 477
rect 270 310 350 326
rect 270 276 300 310
rect 334 276 350 310
rect 270 264 350 276
rect 300 260 350 264
<< polycont >>
rect 60 422 94 456
rect 180 350 214 384
rect 300 276 334 310
<< locali >>
rect 44 422 60 456
rect 94 422 110 456
rect 164 350 180 384
rect 214 350 230 384
rect 164 276 180 310
rect 214 276 300 310
rect 334 276 350 310
<< viali >>
rect 60 422 94 456
rect 180 350 214 384
rect 180 276 214 310
<< metal1 >>
rect 0 615 394 649
rect 48 587 82 615
rect 224 587 258 615
rect 136 475 170 503
rect 312 475 346 503
rect 0 456 106 462
rect 0 428 60 456
rect 48 422 60 428
rect 94 422 106 456
rect 136 441 346 475
rect 48 416 106 422
rect 312 397 346 441
rect 168 384 226 390
rect 0 350 180 384
rect 214 350 226 384
rect 168 344 226 350
rect 312 363 394 397
rect 168 310 226 316
rect 0 276 180 310
rect 214 276 226 310
rect 168 270 226 276
rect 312 238 346 363
rect 48 125 82 154
rect 0 91 394 125
use sky130_fd_pr__nfet_01v8_A6LSUL  m1 ~/Desktop/FabRAM/FE/sram130/common
timestamp 1702396496
transform 1 0 109 0 1 196
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_A6LSUL  m2
timestamp 1702396496
transform 1 0 197 0 1 196
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_A6LSUL  m3
timestamp 1702396496
transform 1 0 285 0 1 196
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_4Y88KP  m4 ~/Desktop/FabRAM/FE/sram130/common
timestamp 1702396496
transform 1 0 109 0 1 545
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m5
timestamp 1702396496
transform -1 0 197 0 1 545
box -109 -104 109 104
use sky130_fd_pr__pfet_01v8_4Y88KP  m6
timestamp 1702396496
transform 1 0 285 0 1 545
box -109 -104 109 104
<< labels >>
rlabel metal1 0 615 34 649 0 VDD
rlabel metal1 0 91 34 125 0 VSS
rlabel metal1 360 363 394 397 0 Y
rlabel metal1 0 350 34 384 0 B
rlabel metal1 0 276 34 310 0 C
rlabel metal1 0 428 34 462 0 A
<< end >>
