magic
tech sky130A
magscale 1 2
timestamp 1702830337
<< nwell >>
rect 0 2369 1345 2577
rect 0 1783 1345 1991
rect 0 1173 1345 1381
rect 0 583 1345 791
<< nmos >>
rect 206 2082 236 2166
rect 803 2082 833 2166
rect 891 2082 921 2166
rect 1221 2082 1251 2166
rect 206 1496 236 1580
rect 803 1496 833 1580
rect 891 1496 921 1580
rect 1221 1496 1251 1580
rect 206 886 236 970
rect 803 886 833 970
rect 891 886 921 970
rect 1221 886 1251 970
rect 206 296 236 380
rect 803 296 833 380
rect 891 296 921 380
rect 1221 296 1251 380
<< pmos >>
rect 206 2431 236 2515
rect 803 2431 833 2515
rect 891 2431 921 2515
rect 1221 2431 1251 2515
rect 206 1845 236 1929
rect 803 1845 833 1929
rect 891 1845 921 1929
rect 1221 1845 1251 1929
rect 206 1235 236 1319
rect 803 1235 833 1319
rect 891 1235 921 1319
rect 1221 1235 1251 1319
rect 206 645 236 729
rect 803 645 833 729
rect 891 645 921 729
rect 1221 645 1251 729
<< ndiff >>
rect 148 2154 206 2166
rect 148 2094 160 2154
rect 194 2094 206 2154
rect 148 2082 206 2094
rect 236 2154 294 2166
rect 236 2094 248 2154
rect 282 2094 294 2154
rect 236 2082 294 2094
rect 745 2154 803 2166
rect 745 2094 757 2154
rect 791 2094 803 2154
rect 745 2082 803 2094
rect 833 2154 891 2166
rect 833 2094 845 2154
rect 879 2094 891 2154
rect 833 2082 891 2094
rect 921 2154 979 2166
rect 921 2094 933 2154
rect 967 2094 979 2154
rect 921 2082 979 2094
rect 1163 2154 1221 2166
rect 1163 2094 1175 2154
rect 1209 2094 1221 2154
rect 1163 2082 1221 2094
rect 1251 2154 1309 2166
rect 1251 2094 1263 2154
rect 1297 2094 1309 2154
rect 1251 2082 1309 2094
rect 148 1568 206 1580
rect 148 1508 160 1568
rect 194 1508 206 1568
rect 148 1496 206 1508
rect 236 1568 294 1580
rect 236 1508 248 1568
rect 282 1508 294 1568
rect 236 1496 294 1508
rect 745 1568 803 1580
rect 745 1508 757 1568
rect 791 1508 803 1568
rect 745 1496 803 1508
rect 833 1568 891 1580
rect 833 1508 845 1568
rect 879 1508 891 1568
rect 833 1496 891 1508
rect 921 1568 979 1580
rect 921 1508 933 1568
rect 967 1508 979 1568
rect 921 1496 979 1508
rect 1163 1568 1221 1580
rect 1163 1508 1175 1568
rect 1209 1508 1221 1568
rect 1163 1496 1221 1508
rect 1251 1568 1309 1580
rect 1251 1508 1263 1568
rect 1297 1508 1309 1568
rect 1251 1496 1309 1508
rect 148 958 206 970
rect 148 898 160 958
rect 194 898 206 958
rect 148 886 206 898
rect 236 958 294 970
rect 236 898 248 958
rect 282 898 294 958
rect 236 886 294 898
rect 745 958 803 970
rect 745 898 757 958
rect 791 898 803 958
rect 745 886 803 898
rect 833 958 891 970
rect 833 898 845 958
rect 879 898 891 958
rect 833 886 891 898
rect 921 958 979 970
rect 921 898 933 958
rect 967 898 979 958
rect 921 886 979 898
rect 1163 958 1221 970
rect 1163 898 1175 958
rect 1209 898 1221 958
rect 1163 886 1221 898
rect 1251 958 1309 970
rect 1251 898 1263 958
rect 1297 898 1309 958
rect 1251 886 1309 898
rect 148 368 206 380
rect 148 308 160 368
rect 194 308 206 368
rect 148 296 206 308
rect 236 368 294 380
rect 236 308 248 368
rect 282 308 294 368
rect 236 296 294 308
rect 745 368 803 380
rect 745 308 757 368
rect 791 308 803 368
rect 745 296 803 308
rect 833 368 891 380
rect 833 308 845 368
rect 879 308 891 368
rect 833 296 891 308
rect 921 368 979 380
rect 921 308 933 368
rect 967 308 979 368
rect 921 296 979 308
rect 1163 368 1221 380
rect 1163 308 1175 368
rect 1209 308 1221 368
rect 1163 296 1221 308
rect 1251 368 1309 380
rect 1251 308 1263 368
rect 1297 308 1309 368
rect 1251 296 1309 308
<< pdiff >>
rect 148 2503 206 2515
rect 148 2443 160 2503
rect 194 2443 206 2503
rect 148 2431 206 2443
rect 236 2503 294 2515
rect 236 2443 248 2503
rect 282 2443 294 2503
rect 236 2431 294 2443
rect 745 2503 803 2515
rect 745 2443 757 2503
rect 791 2443 803 2503
rect 745 2431 803 2443
rect 833 2503 891 2515
rect 833 2443 845 2503
rect 879 2443 891 2503
rect 833 2431 891 2443
rect 921 2503 979 2515
rect 921 2443 933 2503
rect 967 2443 979 2503
rect 921 2431 979 2443
rect 1163 2503 1221 2515
rect 1163 2443 1175 2503
rect 1209 2443 1221 2503
rect 1163 2431 1221 2443
rect 1251 2503 1309 2515
rect 1251 2443 1263 2503
rect 1297 2443 1309 2503
rect 1251 2431 1309 2443
rect 148 1917 206 1929
rect 148 1857 160 1917
rect 194 1857 206 1917
rect 148 1845 206 1857
rect 236 1917 294 1929
rect 236 1857 248 1917
rect 282 1857 294 1917
rect 236 1845 294 1857
rect 745 1917 803 1929
rect 745 1857 757 1917
rect 791 1857 803 1917
rect 745 1845 803 1857
rect 833 1917 891 1929
rect 833 1857 845 1917
rect 879 1857 891 1917
rect 833 1845 891 1857
rect 921 1917 979 1929
rect 921 1857 933 1917
rect 967 1857 979 1917
rect 921 1845 979 1857
rect 1163 1917 1221 1929
rect 1163 1857 1175 1917
rect 1209 1857 1221 1917
rect 1163 1845 1221 1857
rect 1251 1917 1309 1929
rect 1251 1857 1263 1917
rect 1297 1857 1309 1917
rect 1251 1845 1309 1857
rect 148 1307 206 1319
rect 148 1247 160 1307
rect 194 1247 206 1307
rect 148 1235 206 1247
rect 236 1307 294 1319
rect 236 1247 248 1307
rect 282 1247 294 1307
rect 236 1235 294 1247
rect 745 1307 803 1319
rect 745 1247 757 1307
rect 791 1247 803 1307
rect 745 1235 803 1247
rect 833 1307 891 1319
rect 833 1247 845 1307
rect 879 1247 891 1307
rect 833 1235 891 1247
rect 921 1307 979 1319
rect 921 1247 933 1307
rect 967 1247 979 1307
rect 921 1235 979 1247
rect 1163 1307 1221 1319
rect 1163 1247 1175 1307
rect 1209 1247 1221 1307
rect 1163 1235 1221 1247
rect 1251 1307 1309 1319
rect 1251 1247 1263 1307
rect 1297 1247 1309 1307
rect 1251 1235 1309 1247
rect 148 717 206 729
rect 148 657 160 717
rect 194 657 206 717
rect 148 645 206 657
rect 236 717 294 729
rect 236 657 248 717
rect 282 657 294 717
rect 236 645 294 657
rect 745 717 803 729
rect 745 657 757 717
rect 791 657 803 717
rect 745 645 803 657
rect 833 717 891 729
rect 833 657 845 717
rect 879 657 891 717
rect 833 645 891 657
rect 921 717 979 729
rect 921 657 933 717
rect 967 657 979 717
rect 921 645 979 657
rect 1163 717 1221 729
rect 1163 657 1175 717
rect 1209 657 1221 717
rect 1163 645 1221 657
rect 1251 717 1309 729
rect 1251 657 1263 717
rect 1297 657 1309 717
rect 1251 645 1309 657
<< ndiffc >>
rect 160 2094 194 2154
rect 248 2094 282 2154
rect 757 2094 791 2154
rect 845 2094 879 2154
rect 933 2094 967 2154
rect 1175 2094 1209 2154
rect 1263 2094 1297 2154
rect 160 1508 194 1568
rect 248 1508 282 1568
rect 757 1508 791 1568
rect 845 1508 879 1568
rect 933 1508 967 1568
rect 1175 1508 1209 1568
rect 1263 1508 1297 1568
rect 160 898 194 958
rect 248 898 282 958
rect 757 898 791 958
rect 845 898 879 958
rect 933 898 967 958
rect 1175 898 1209 958
rect 1263 898 1297 958
rect 160 308 194 368
rect 248 308 282 368
rect 757 308 791 368
rect 845 308 879 368
rect 933 308 967 368
rect 1175 308 1209 368
rect 1263 308 1297 368
<< pdiffc >>
rect 160 2443 194 2503
rect 248 2443 282 2503
rect 757 2443 791 2503
rect 845 2443 879 2503
rect 933 2443 967 2503
rect 1175 2443 1209 2503
rect 1263 2443 1297 2503
rect 160 1857 194 1917
rect 248 1857 282 1917
rect 757 1857 791 1917
rect 845 1857 879 1917
rect 933 1857 967 1917
rect 1175 1857 1209 1917
rect 1263 1857 1297 1917
rect 160 1247 194 1307
rect 248 1247 282 1307
rect 757 1247 791 1307
rect 845 1247 879 1307
rect 933 1247 967 1307
rect 1175 1247 1209 1307
rect 1263 1247 1297 1307
rect 160 657 194 717
rect 248 657 282 717
rect 757 657 791 717
rect 845 657 879 717
rect 933 657 967 717
rect 1175 657 1209 717
rect 1263 657 1297 717
<< psubdiff >>
rect 36 2154 94 2178
rect 36 2094 48 2154
rect 82 2094 94 2154
rect 36 2070 94 2094
rect 1051 2154 1109 2178
rect 1051 2094 1063 2154
rect 1097 2094 1109 2154
rect 1051 2070 1109 2094
rect 36 1568 94 1592
rect 36 1508 48 1568
rect 82 1508 94 1568
rect 36 1484 94 1508
rect 1051 1568 1109 1592
rect 1051 1508 1063 1568
rect 1097 1508 1109 1568
rect 1051 1484 1109 1508
rect 36 958 94 982
rect 36 898 48 958
rect 82 898 94 958
rect 36 874 94 898
rect 1051 958 1109 982
rect 1051 898 1063 958
rect 1097 898 1109 958
rect 1051 874 1109 898
rect 36 368 94 392
rect 36 308 48 368
rect 82 308 94 368
rect 36 284 94 308
rect 1051 368 1109 392
rect 1051 308 1063 368
rect 1097 308 1109 368
rect 1051 284 1109 308
<< nsubdiff >>
rect 36 2503 94 2527
rect 36 2443 48 2503
rect 82 2443 94 2503
rect 36 2419 94 2443
rect 1051 2503 1109 2527
rect 1051 2443 1063 2503
rect 1097 2443 1109 2503
rect 1051 2419 1109 2443
rect 36 1917 94 1941
rect 36 1857 48 1917
rect 82 1857 94 1917
rect 36 1833 94 1857
rect 1051 1917 1109 1941
rect 1051 1857 1063 1917
rect 1097 1857 1109 1917
rect 1051 1833 1109 1857
rect 36 1307 94 1331
rect 36 1247 48 1307
rect 82 1247 94 1307
rect 36 1223 94 1247
rect 1051 1307 1109 1331
rect 1051 1247 1063 1307
rect 1097 1247 1109 1307
rect 1051 1223 1109 1247
rect 36 717 94 741
rect 36 657 48 717
rect 82 657 94 717
rect 36 633 94 657
rect 1051 717 1109 741
rect 1051 657 1063 717
rect 1097 657 1109 717
rect 1051 633 1109 657
<< psubdiffcont >>
rect 48 2094 82 2154
rect 1063 2094 1097 2154
rect 48 1508 82 1568
rect 1063 1508 1097 1568
rect 48 898 82 958
rect 1063 898 1097 958
rect 48 308 82 368
rect 1063 308 1097 368
<< nsubdiffcont >>
rect 48 2443 82 2503
rect 1063 2443 1097 2503
rect 48 1857 82 1917
rect 1063 1857 1097 1917
rect 48 1247 82 1307
rect 1063 1247 1097 1307
rect 48 657 82 717
rect 1063 657 1097 717
<< poly >>
rect 206 2515 236 2541
rect 803 2515 833 2541
rect 891 2515 921 2541
rect 1221 2515 1251 2541
rect 206 2341 236 2431
rect 803 2399 833 2431
rect 145 2325 236 2341
rect 753 2383 833 2399
rect 753 2349 769 2383
rect 803 2349 833 2383
rect 753 2333 833 2349
rect 145 2291 161 2325
rect 195 2291 236 2325
rect 145 2275 236 2291
rect 206 2166 236 2275
rect 803 2166 833 2333
rect 891 2254 921 2431
rect 1221 2341 1251 2431
rect 1160 2325 1251 2341
rect 1160 2291 1176 2325
rect 1210 2291 1251 2325
rect 1160 2275 1251 2291
rect 891 2238 971 2254
rect 891 2204 921 2238
rect 955 2204 971 2238
rect 891 2188 971 2204
rect 891 2166 921 2188
rect 1221 2166 1251 2275
rect 206 2056 236 2082
rect 803 2056 833 2082
rect 891 2056 921 2082
rect 1221 2056 1251 2082
rect 206 1929 236 1955
rect 803 1929 833 1955
rect 891 1929 921 1955
rect 1221 1929 1251 1955
rect 206 1755 236 1845
rect 803 1813 833 1845
rect 145 1739 236 1755
rect 753 1797 833 1813
rect 753 1763 769 1797
rect 803 1763 833 1797
rect 753 1747 833 1763
rect 145 1705 161 1739
rect 195 1705 236 1739
rect 145 1689 236 1705
rect 206 1580 236 1689
rect 803 1580 833 1747
rect 891 1668 921 1845
rect 1221 1755 1251 1845
rect 1160 1739 1251 1755
rect 1160 1705 1176 1739
rect 1210 1705 1251 1739
rect 1160 1689 1251 1705
rect 891 1652 971 1668
rect 891 1618 921 1652
rect 955 1618 971 1652
rect 891 1602 971 1618
rect 891 1580 921 1602
rect 1221 1580 1251 1689
rect 206 1470 236 1496
rect 803 1470 833 1496
rect 891 1470 921 1496
rect 1221 1470 1251 1496
rect 206 1319 236 1345
rect 803 1319 833 1345
rect 891 1319 921 1345
rect 1221 1319 1251 1345
rect 206 1145 236 1235
rect 803 1203 833 1235
rect 145 1129 236 1145
rect 753 1187 833 1203
rect 753 1153 769 1187
rect 803 1153 833 1187
rect 753 1137 833 1153
rect 145 1095 161 1129
rect 195 1095 236 1129
rect 145 1079 236 1095
rect 206 970 236 1079
rect 803 970 833 1137
rect 891 1058 921 1235
rect 1221 1145 1251 1235
rect 1160 1129 1251 1145
rect 1160 1095 1176 1129
rect 1210 1095 1251 1129
rect 1160 1079 1251 1095
rect 891 1042 971 1058
rect 891 1008 921 1042
rect 955 1008 971 1042
rect 891 992 971 1008
rect 891 970 921 992
rect 1221 970 1251 1079
rect 206 860 236 886
rect 803 860 833 886
rect 891 860 921 886
rect 1221 860 1251 886
rect 206 729 236 755
rect 803 729 833 755
rect 891 729 921 755
rect 1221 729 1251 755
rect 206 555 236 645
rect 803 613 833 645
rect 145 539 236 555
rect 753 597 833 613
rect 753 563 769 597
rect 803 563 833 597
rect 753 547 833 563
rect 145 505 161 539
rect 195 505 236 539
rect 145 489 236 505
rect 206 380 236 489
rect 803 380 833 547
rect 891 468 921 645
rect 1221 555 1251 645
rect 1160 539 1251 555
rect 1160 505 1176 539
rect 1210 505 1251 539
rect 1160 489 1251 505
rect 891 452 971 468
rect 891 418 921 452
rect 955 418 971 452
rect 891 402 971 418
rect 891 380 921 402
rect 1221 380 1251 489
rect 206 270 236 296
rect 803 270 833 296
rect 891 270 921 296
rect 1221 270 1251 296
<< polycont >>
rect 769 2349 803 2383
rect 161 2291 195 2325
rect 1176 2291 1210 2325
rect 921 2204 955 2238
rect 769 1763 803 1797
rect 161 1705 195 1739
rect 1176 1705 1210 1739
rect 921 1618 955 1652
rect 769 1153 803 1187
rect 161 1095 195 1129
rect 1176 1095 1210 1129
rect 921 1008 955 1042
rect 769 563 803 597
rect 161 505 195 539
rect 1176 505 1210 539
rect 921 418 955 452
<< locali >>
rect 36 2503 194 2519
rect 36 2443 48 2503
rect 82 2443 160 2503
rect 36 2427 194 2443
rect 248 2503 282 2519
rect 248 2325 282 2443
rect 757 2503 791 2519
rect 757 2427 791 2443
rect 845 2503 879 2519
rect 845 2427 879 2443
rect 933 2503 967 2519
rect 933 2427 967 2443
rect 1051 2503 1209 2519
rect 1051 2443 1063 2503
rect 1097 2443 1175 2503
rect 1051 2427 1209 2443
rect 1263 2503 1297 2519
rect 753 2349 769 2383
rect 803 2349 819 2383
rect 1263 2325 1297 2443
rect 145 2291 161 2325
rect 195 2291 211 2325
rect 1160 2291 1176 2325
rect 1210 2291 1226 2325
rect 48 2154 194 2170
rect 82 2094 160 2154
rect 48 2078 194 2094
rect 248 2154 282 2291
rect 757 2204 769 2238
rect 803 2204 921 2238
rect 955 2204 971 2238
rect 248 2078 282 2094
rect 757 2154 791 2170
rect 757 2078 791 2094
rect 845 2154 879 2170
rect 845 2078 879 2094
rect 933 2154 967 2170
rect 933 2078 967 2094
rect 1063 2154 1209 2170
rect 1097 2094 1175 2154
rect 1063 2078 1209 2094
rect 1263 2154 1297 2291
rect 1263 2078 1297 2094
rect 36 1917 194 1933
rect 36 1857 48 1917
rect 82 1857 160 1917
rect 36 1841 194 1857
rect 248 1917 282 1933
rect 248 1739 282 1857
rect 757 1917 791 1933
rect 757 1841 791 1857
rect 845 1917 879 1933
rect 845 1841 879 1857
rect 933 1917 967 1933
rect 933 1841 967 1857
rect 1051 1917 1209 1933
rect 1051 1857 1063 1917
rect 1097 1857 1175 1917
rect 1051 1841 1209 1857
rect 1263 1917 1297 1933
rect 753 1763 769 1797
rect 803 1763 819 1797
rect 1263 1739 1297 1857
rect 145 1705 161 1739
rect 195 1705 211 1739
rect 1160 1705 1176 1739
rect 1210 1705 1226 1739
rect 48 1568 194 1584
rect 82 1508 160 1568
rect 48 1492 194 1508
rect 248 1568 282 1705
rect 757 1618 769 1652
rect 803 1618 921 1652
rect 955 1618 971 1652
rect 248 1492 282 1508
rect 757 1568 791 1584
rect 757 1492 791 1508
rect 845 1568 879 1584
rect 845 1492 879 1508
rect 933 1568 967 1584
rect 933 1492 967 1508
rect 1063 1568 1209 1584
rect 1097 1508 1175 1568
rect 1063 1492 1209 1508
rect 1263 1568 1297 1705
rect 1263 1492 1297 1508
rect 36 1307 194 1323
rect 36 1247 48 1307
rect 82 1247 160 1307
rect 36 1231 194 1247
rect 248 1307 282 1323
rect 248 1129 282 1247
rect 757 1307 791 1323
rect 757 1231 791 1247
rect 845 1307 879 1323
rect 845 1231 879 1247
rect 933 1307 967 1323
rect 933 1231 967 1247
rect 1051 1307 1209 1323
rect 1051 1247 1063 1307
rect 1097 1247 1175 1307
rect 1051 1231 1209 1247
rect 1263 1307 1297 1323
rect 753 1153 769 1187
rect 803 1153 819 1187
rect 1263 1129 1297 1247
rect 145 1095 161 1129
rect 195 1095 211 1129
rect 1160 1095 1176 1129
rect 1210 1095 1226 1129
rect 48 958 194 974
rect 82 898 160 958
rect 48 882 194 898
rect 248 958 282 1095
rect 757 1008 769 1042
rect 803 1008 921 1042
rect 955 1008 971 1042
rect 248 882 282 898
rect 757 958 791 974
rect 757 882 791 898
rect 845 958 879 974
rect 845 882 879 898
rect 933 958 967 974
rect 933 882 967 898
rect 1063 958 1209 974
rect 1097 898 1175 958
rect 1063 882 1209 898
rect 1263 958 1297 1095
rect 1263 882 1297 898
rect 36 717 194 733
rect 36 657 48 717
rect 82 657 160 717
rect 36 641 194 657
rect 248 717 282 733
rect 248 539 282 657
rect 757 717 791 733
rect 757 641 791 657
rect 845 717 879 733
rect 845 641 879 657
rect 933 717 967 733
rect 933 641 967 657
rect 1051 717 1209 733
rect 1051 657 1063 717
rect 1097 657 1175 717
rect 1051 641 1209 657
rect 1263 717 1297 733
rect 753 563 769 597
rect 803 563 819 597
rect 1263 539 1297 657
rect 145 505 161 539
rect 195 505 211 539
rect 1160 505 1176 539
rect 1210 505 1226 539
rect 48 368 194 384
rect 82 308 160 368
rect 48 292 194 308
rect 248 368 282 505
rect 757 418 769 452
rect 803 418 921 452
rect 955 418 971 452
rect 248 292 282 308
rect 757 368 791 384
rect 757 292 791 308
rect 845 368 879 384
rect 845 292 879 308
rect 933 368 967 384
rect 933 292 967 308
rect 1063 368 1209 384
rect 1097 308 1175 368
rect 1063 292 1209 308
rect 1263 368 1297 505
rect 1263 292 1297 308
<< viali >>
rect 160 2443 194 2503
rect 248 2443 282 2503
rect 757 2443 791 2503
rect 845 2443 879 2503
rect 933 2443 967 2503
rect 1175 2443 1209 2503
rect 1263 2443 1297 2503
rect 769 2349 803 2383
rect 161 2291 195 2325
rect 248 2291 282 2325
rect 1176 2291 1210 2325
rect 1263 2291 1297 2325
rect 160 2094 194 2154
rect 769 2204 803 2238
rect 248 2094 282 2154
rect 757 2094 791 2154
rect 845 2094 879 2154
rect 933 2094 967 2154
rect 1175 2094 1209 2154
rect 1263 2094 1297 2154
rect 160 1857 194 1917
rect 248 1857 282 1917
rect 757 1857 791 1917
rect 845 1857 879 1917
rect 933 1857 967 1917
rect 1175 1857 1209 1917
rect 1263 1857 1297 1917
rect 769 1763 803 1797
rect 161 1705 195 1739
rect 248 1705 282 1739
rect 1176 1705 1210 1739
rect 1263 1705 1297 1739
rect 160 1508 194 1568
rect 769 1618 803 1652
rect 248 1508 282 1568
rect 757 1508 791 1568
rect 845 1508 879 1568
rect 933 1508 967 1568
rect 1175 1508 1209 1568
rect 1263 1508 1297 1568
rect 160 1247 194 1307
rect 248 1247 282 1307
rect 757 1247 791 1307
rect 845 1247 879 1307
rect 933 1247 967 1307
rect 1175 1247 1209 1307
rect 1263 1247 1297 1307
rect 769 1153 803 1187
rect 161 1095 195 1129
rect 248 1095 282 1129
rect 1176 1095 1210 1129
rect 1263 1095 1297 1129
rect 160 898 194 958
rect 769 1008 803 1042
rect 248 898 282 958
rect 757 898 791 958
rect 845 898 879 958
rect 933 898 967 958
rect 1175 898 1209 958
rect 1263 898 1297 958
rect 160 657 194 717
rect 248 657 282 717
rect 757 657 791 717
rect 845 657 879 717
rect 933 657 967 717
rect 1175 657 1209 717
rect 1263 657 1297 717
rect 769 563 803 597
rect 161 505 195 539
rect 248 505 282 539
rect 1176 505 1210 539
rect 1263 505 1297 539
rect 160 308 194 368
rect 769 418 803 452
rect 248 308 282 368
rect 757 308 791 368
rect 845 308 879 368
rect 933 308 967 368
rect 1175 308 1209 368
rect 1263 308 1297 368
<< metal1 >>
rect 0 2543 647 2577
rect 160 2515 194 2543
rect 637 2525 647 2543
rect 699 2543 1345 2577
rect 699 2525 709 2543
rect 757 2515 791 2543
rect 933 2515 967 2543
rect 1175 2515 1209 2543
rect 154 2503 200 2515
rect 154 2443 160 2503
rect 194 2443 200 2503
rect 154 2431 200 2443
rect 242 2503 288 2515
rect 242 2443 248 2503
rect 282 2443 288 2503
rect 242 2431 288 2443
rect 751 2503 797 2515
rect 751 2443 757 2503
rect 791 2443 797 2503
rect 751 2431 797 2443
rect 839 2503 885 2515
rect 839 2443 845 2503
rect 879 2443 885 2503
rect 839 2431 885 2443
rect 927 2503 973 2515
rect 927 2443 933 2503
rect 967 2443 973 2503
rect 927 2431 973 2443
rect 1169 2503 1215 2515
rect 1169 2443 1175 2503
rect 1209 2443 1215 2503
rect 1169 2431 1215 2443
rect 1257 2503 1303 2515
rect 1257 2443 1263 2503
rect 1297 2443 1303 2503
rect 1257 2431 1303 2443
rect 477 2349 487 2401
rect 539 2383 549 2401
rect 757 2383 815 2389
rect 539 2349 769 2383
rect 803 2349 815 2383
rect 757 2343 815 2349
rect 272 2331 282 2334
rect 149 2325 207 2331
rect 0 2291 161 2325
rect 195 2291 207 2325
rect 149 2285 207 2291
rect 236 2325 282 2331
rect 236 2291 248 2325
rect 236 2285 282 2291
rect 272 2282 282 2285
rect 334 2282 344 2334
rect 845 2325 879 2431
rect 1299 2331 1309 2334
rect 1164 2325 1222 2331
rect 845 2291 1176 2325
rect 1210 2291 1222 2325
rect 397 2204 407 2256
rect 459 2238 469 2256
rect 757 2238 815 2244
rect 459 2204 769 2238
rect 803 2204 815 2238
rect 757 2198 815 2204
rect 933 2166 967 2291
rect 1164 2285 1222 2291
rect 1251 2325 1309 2331
rect 1251 2291 1263 2325
rect 1297 2291 1309 2325
rect 1251 2285 1309 2291
rect 1299 2282 1309 2285
rect 1361 2282 1371 2334
rect 154 2154 200 2166
rect 154 2094 160 2154
rect 194 2094 200 2154
rect 154 2082 200 2094
rect 242 2154 288 2166
rect 242 2094 248 2154
rect 282 2094 288 2154
rect 242 2082 288 2094
rect 751 2154 797 2166
rect 751 2094 757 2154
rect 791 2094 797 2154
rect 751 2082 797 2094
rect 839 2154 885 2166
rect 839 2094 845 2154
rect 879 2094 885 2154
rect 839 2082 885 2094
rect 927 2154 973 2166
rect 927 2094 933 2154
rect 967 2094 973 2154
rect 927 2082 973 2094
rect 1169 2154 1215 2166
rect 1169 2094 1175 2154
rect 1209 2094 1215 2154
rect 1169 2082 1215 2094
rect 1257 2154 1303 2166
rect 1257 2094 1263 2154
rect 1297 2094 1303 2154
rect 1257 2082 1303 2094
rect 160 2053 194 2082
rect 557 2053 567 2071
rect 0 2019 567 2053
rect 619 2053 629 2071
rect 757 2053 791 2082
rect 1175 2053 1209 2082
rect 619 2019 1345 2053
rect 0 1957 647 1991
rect 160 1929 194 1957
rect 637 1939 647 1957
rect 699 1957 1345 1991
rect 699 1939 709 1957
rect 757 1929 791 1957
rect 933 1929 967 1957
rect 1175 1929 1209 1957
rect 154 1917 200 1929
rect 154 1857 160 1917
rect 194 1857 200 1917
rect 154 1845 200 1857
rect 242 1917 288 1929
rect 242 1857 248 1917
rect 282 1857 288 1917
rect 242 1845 288 1857
rect 751 1917 797 1929
rect 751 1857 757 1917
rect 791 1857 797 1917
rect 751 1845 797 1857
rect 839 1917 885 1929
rect 839 1857 845 1917
rect 879 1857 885 1917
rect 839 1845 885 1857
rect 927 1917 973 1929
rect 927 1857 933 1917
rect 967 1857 973 1917
rect 927 1845 973 1857
rect 1169 1917 1215 1929
rect 1169 1857 1175 1917
rect 1209 1857 1215 1917
rect 1169 1845 1215 1857
rect 1257 1917 1303 1929
rect 1257 1857 1263 1917
rect 1297 1857 1303 1917
rect 1257 1845 1303 1857
rect 477 1763 487 1815
rect 539 1797 549 1815
rect 757 1797 815 1803
rect 539 1763 769 1797
rect 803 1763 815 1797
rect 149 1739 207 1745
rect 0 1705 161 1739
rect 195 1705 207 1739
rect 149 1699 207 1705
rect 236 1739 294 1745
rect 477 1739 505 1763
rect 757 1757 815 1763
rect 236 1705 248 1739
rect 282 1705 505 1739
rect 845 1739 879 1845
rect 1299 1745 1309 1748
rect 1164 1739 1222 1745
rect 845 1705 1176 1739
rect 1210 1705 1222 1739
rect 236 1699 294 1705
rect 161 1662 195 1699
rect 477 1662 487 1671
rect 161 1628 487 1662
rect 477 1619 487 1628
rect 539 1619 549 1671
rect 757 1652 815 1658
rect 647 1618 769 1652
rect 803 1618 815 1652
rect 154 1568 200 1580
rect 154 1508 160 1568
rect 194 1508 200 1568
rect 154 1496 200 1508
rect 242 1568 288 1580
rect 242 1508 248 1568
rect 282 1508 288 1568
rect 317 1533 327 1585
rect 379 1567 389 1585
rect 647 1567 681 1618
rect 757 1612 815 1618
rect 933 1580 967 1705
rect 1164 1699 1222 1705
rect 1251 1739 1309 1745
rect 1251 1705 1263 1739
rect 1297 1705 1309 1739
rect 1251 1699 1309 1705
rect 1299 1696 1309 1699
rect 1361 1696 1371 1748
rect 379 1533 681 1567
rect 751 1568 797 1580
rect 242 1496 288 1508
rect 751 1508 757 1568
rect 791 1508 797 1568
rect 751 1496 797 1508
rect 839 1568 885 1580
rect 839 1508 845 1568
rect 879 1508 885 1568
rect 839 1496 885 1508
rect 927 1568 973 1580
rect 927 1508 933 1568
rect 967 1508 973 1568
rect 927 1496 973 1508
rect 1169 1568 1215 1580
rect 1169 1508 1175 1568
rect 1209 1508 1215 1568
rect 1169 1496 1215 1508
rect 1257 1568 1303 1580
rect 1257 1508 1263 1568
rect 1297 1508 1303 1568
rect 1257 1496 1303 1508
rect 160 1467 194 1496
rect 557 1467 567 1495
rect 0 1443 567 1467
rect 619 1467 629 1495
rect 757 1467 791 1496
rect 1175 1467 1209 1496
rect 619 1443 1345 1467
rect 0 1433 1345 1443
rect 327 1432 455 1433
rect 0 1347 647 1381
rect 160 1319 194 1347
rect 637 1329 647 1347
rect 699 1347 1345 1381
rect 699 1329 709 1347
rect 757 1319 791 1347
rect 933 1319 967 1347
rect 1175 1319 1209 1347
rect 154 1307 200 1319
rect 154 1247 160 1307
rect 194 1247 200 1307
rect 154 1235 200 1247
rect 242 1307 288 1319
rect 242 1247 248 1307
rect 282 1247 288 1307
rect 242 1235 288 1247
rect 751 1307 797 1319
rect 751 1247 757 1307
rect 791 1247 797 1307
rect 751 1235 797 1247
rect 839 1307 885 1319
rect 839 1247 845 1307
rect 879 1247 885 1307
rect 839 1235 885 1247
rect 927 1307 973 1319
rect 927 1247 933 1307
rect 967 1247 973 1307
rect 927 1235 973 1247
rect 1169 1307 1215 1319
rect 1169 1247 1175 1307
rect 1209 1247 1215 1307
rect 1169 1235 1215 1247
rect 1257 1307 1303 1319
rect 1257 1247 1263 1307
rect 1297 1247 1303 1307
rect 1257 1235 1303 1247
rect 477 1153 487 1205
rect 539 1187 549 1205
rect 757 1187 815 1193
rect 539 1153 769 1187
rect 803 1153 815 1187
rect 757 1147 815 1153
rect 149 1129 207 1135
rect 0 1095 161 1129
rect 195 1095 207 1129
rect 149 1089 207 1095
rect 236 1129 294 1135
rect 845 1129 879 1235
rect 1299 1135 1309 1138
rect 1164 1129 1222 1135
rect 236 1095 248 1129
rect 282 1095 431 1129
rect 845 1095 1176 1129
rect 1210 1095 1222 1129
rect 236 1089 294 1095
rect 161 1034 195 1089
rect 397 1060 431 1095
rect 161 1000 351 1034
rect 397 1008 407 1060
rect 459 1042 469 1060
rect 757 1042 815 1048
rect 459 1008 769 1042
rect 803 1008 815 1042
rect 757 1002 815 1008
rect 154 958 200 970
rect 154 898 160 958
rect 194 898 200 958
rect 154 886 200 898
rect 242 958 288 970
rect 242 898 248 958
rect 282 898 288 958
rect 317 957 351 1000
rect 933 970 967 1095
rect 1164 1089 1222 1095
rect 1251 1129 1309 1135
rect 1251 1095 1263 1129
rect 1297 1095 1309 1129
rect 1251 1089 1309 1095
rect 1299 1086 1309 1089
rect 1361 1086 1371 1138
rect 751 958 797 970
rect 317 905 327 957
rect 379 905 389 957
rect 242 886 288 898
rect 751 898 757 958
rect 791 898 797 958
rect 751 886 797 898
rect 839 958 885 970
rect 839 898 845 958
rect 879 898 885 958
rect 839 886 885 898
rect 927 958 973 970
rect 927 898 933 958
rect 967 898 973 958
rect 927 886 973 898
rect 1169 958 1215 970
rect 1169 898 1175 958
rect 1209 898 1215 958
rect 1169 886 1215 898
rect 1257 958 1303 970
rect 1257 898 1263 958
rect 1297 898 1303 958
rect 1257 886 1303 898
rect 160 857 194 886
rect 557 857 567 885
rect 0 833 567 857
rect 619 857 629 885
rect 757 857 791 886
rect 1175 857 1209 886
rect 619 833 1345 857
rect 0 823 1345 833
rect 160 757 647 791
rect 160 729 194 757
rect 637 739 647 757
rect 699 757 1345 791
rect 699 739 709 757
rect 757 729 791 757
rect 933 729 967 757
rect 1175 729 1209 757
rect 154 717 200 729
rect 154 657 160 717
rect 194 657 200 717
rect 154 645 200 657
rect 242 717 288 729
rect 242 657 248 717
rect 282 657 288 717
rect 242 645 288 657
rect 751 717 797 729
rect 751 657 757 717
rect 791 657 797 717
rect 751 645 797 657
rect 839 717 885 729
rect 839 657 845 717
rect 879 657 885 717
rect 839 645 885 657
rect 927 717 973 729
rect 927 657 933 717
rect 967 657 973 717
rect 927 645 973 657
rect 1169 717 1215 729
rect 1169 657 1175 717
rect 1209 657 1215 717
rect 1169 645 1215 657
rect 1257 717 1303 729
rect 1257 657 1263 717
rect 1297 657 1303 717
rect 1257 645 1303 657
rect 477 563 487 615
rect 539 597 549 615
rect 757 597 815 603
rect 539 563 769 597
rect 803 563 815 597
rect 757 557 815 563
rect 135 496 145 548
rect 197 496 207 548
rect 236 498 246 550
rect 298 498 330 550
rect 845 539 879 645
rect 1299 545 1309 548
rect 1164 539 1222 545
rect 845 505 1176 539
rect 1210 505 1222 539
rect 316 418 326 470
rect 378 452 388 470
rect 757 452 815 458
rect 378 418 769 452
rect 803 418 815 452
rect 757 412 815 418
rect 933 380 967 505
rect 1164 499 1222 505
rect 1251 539 1309 545
rect 1251 505 1263 539
rect 1297 505 1309 539
rect 1251 499 1309 505
rect 1299 496 1309 499
rect 1361 496 1371 548
rect 154 368 200 380
rect 154 308 160 368
rect 194 308 200 368
rect 154 296 200 308
rect 242 368 288 380
rect 242 308 248 368
rect 282 308 288 368
rect 242 296 288 308
rect 751 368 797 380
rect 751 308 757 368
rect 791 308 797 368
rect 751 296 797 308
rect 839 368 885 380
rect 839 308 845 368
rect 879 308 885 368
rect 839 296 885 308
rect 927 368 973 380
rect 927 308 933 368
rect 967 308 973 368
rect 927 296 973 308
rect 1169 368 1215 380
rect 1169 308 1175 368
rect 1209 308 1215 368
rect 1169 296 1215 308
rect 1257 368 1303 380
rect 1257 308 1263 368
rect 1297 308 1303 368
rect 1257 296 1303 308
rect 160 267 194 296
rect 557 267 567 285
rect 160 233 567 267
rect 619 267 629 285
rect 757 267 791 296
rect 1175 267 1209 296
rect 619 233 1345 267
<< via1 >>
rect 647 2525 699 2577
rect 487 2349 539 2401
rect 282 2282 334 2334
rect 407 2204 459 2256
rect 1309 2282 1361 2334
rect 567 2019 619 2071
rect 647 1939 699 1991
rect 487 1763 539 1815
rect 487 1619 539 1671
rect 327 1533 379 1585
rect 1309 1696 1361 1748
rect 567 1443 619 1495
rect 647 1329 699 1381
rect 487 1153 539 1205
rect 407 1008 459 1060
rect 1309 1086 1361 1138
rect 327 905 379 957
rect 567 833 619 885
rect 647 739 699 791
rect 487 563 539 615
rect 145 539 197 548
rect 145 505 161 539
rect 161 505 195 539
rect 195 505 197 539
rect 145 496 197 505
rect 246 539 298 550
rect 246 505 248 539
rect 248 505 282 539
rect 282 505 298 539
rect 246 498 298 505
rect 326 418 378 470
rect 1309 496 1361 548
rect 567 233 619 285
<< metal2 >>
rect 487 2401 539 2411
rect 282 2334 334 2344
rect 282 1741 334 2282
rect 145 1689 334 1741
rect 407 2256 459 2266
rect 145 548 197 1689
rect 327 1585 379 1595
rect 327 957 379 1533
rect 407 1060 459 2204
rect 487 1815 539 2349
rect 487 1757 539 1763
rect 567 2071 619 2645
rect 407 1000 459 1008
rect 487 1671 539 1679
rect 487 1205 539 1619
rect 145 202 197 496
rect 246 550 298 560
rect 142 192 200 202
rect 142 127 200 136
rect 246 75 298 498
rect 327 480 379 905
rect 487 615 539 1153
rect 487 554 539 563
rect 567 1495 619 2019
rect 567 885 619 1443
rect 326 470 379 480
rect 378 418 379 470
rect 326 408 379 418
rect 567 285 619 833
rect 243 66 301 75
rect 243 0 301 10
rect 567 0 619 233
rect 647 2577 699 2645
rect 647 1991 699 2525
rect 1307 2336 1363 2346
rect 1307 2270 1363 2280
rect 647 1381 699 1939
rect 1307 1750 1363 1760
rect 1307 1684 1363 1694
rect 647 791 699 1329
rect 1307 1140 1363 1150
rect 1307 1074 1363 1084
rect 647 0 699 739
rect 1307 550 1363 560
rect 1307 484 1363 494
<< via2 >>
rect 142 136 200 192
rect 243 10 301 66
rect 1307 2334 1363 2336
rect 1307 2282 1309 2334
rect 1309 2282 1361 2334
rect 1361 2282 1363 2334
rect 1307 2280 1363 2282
rect 1307 1748 1363 1750
rect 1307 1696 1309 1748
rect 1309 1696 1361 1748
rect 1361 1696 1363 1748
rect 1307 1694 1363 1696
rect 1307 1138 1363 1140
rect 1307 1086 1309 1138
rect 1309 1086 1361 1138
rect 1361 1086 1363 1138
rect 1307 1084 1363 1086
rect 1307 548 1363 550
rect 1307 496 1309 548
rect 1309 496 1361 548
rect 1361 496 1363 548
rect 1307 494 1363 496
<< metal3 >>
rect 1297 2336 1462 2341
rect 1297 2280 1307 2336
rect 1363 2280 1462 2336
rect 1297 2275 1462 2280
rect 1297 1750 1462 1755
rect 1297 1694 1307 1750
rect 1363 1694 1462 1750
rect 1297 1689 1462 1694
rect 1297 1140 1462 1145
rect 1297 1084 1307 1140
rect 1363 1084 1462 1140
rect 1297 1079 1462 1084
rect 1297 550 1462 555
rect 1297 494 1307 550
rect 1363 494 1462 550
rect 1297 489 1462 494
rect 132 192 1462 197
rect 132 136 142 192
rect 200 136 1462 192
rect 132 131 1462 136
rect 233 66 1462 71
rect 233 10 243 66
rect 301 10 1462 66
rect 233 5 1462 10
<< labels >>
rlabel metal2 647 2593 699 2645 0 VDD
rlabel metal2 567 2593 619 2645 0 VSS
rlabel metal1 0 2291 34 2325 0 A2
rlabel metal1 0 1705 34 1739 0 A1
rlabel metal1 0 1095 34 1129 0 A0
rlabel metal3 1396 2275 1462 2341 0 Y0
rlabel metal3 1396 1689 1462 1755 0 Y1
rlabel metal3 1396 1079 1462 1145 0 Y2
rlabel metal3 1396 489 1462 555 0 Y3
rlabel metal3 1396 131 1462 197 0 Y4
rlabel metal3 1396 5 1462 71 0 Y5
<< end >>
