magic
tech sky130A
magscale 1 2
timestamp 1703586424
<< nwell >>
rect 0 488 330 696
<< pwell >>
rect 10 311 120 323
rect 10 175 320 311
rect 10 163 120 175
<< nmos >>
rect 206 201 236 285
<< pmos >>
rect 206 550 236 634
<< ndiff >>
rect 148 260 206 285
rect 148 226 160 260
rect 194 226 206 260
rect 148 201 206 226
rect 236 260 294 285
rect 236 226 248 260
rect 282 226 294 260
rect 236 201 294 226
<< pdiff >>
rect 148 609 206 634
rect 148 575 160 609
rect 194 575 206 609
rect 148 550 206 575
rect 236 609 294 634
rect 236 575 248 609
rect 282 575 294 609
rect 236 550 294 575
<< ndiffc >>
rect 160 226 194 260
rect 248 226 282 260
<< pdiffc >>
rect 160 575 194 609
rect 248 575 282 609
<< psubdiff >>
rect 36 260 94 297
rect 36 226 48 260
rect 82 226 94 260
rect 36 189 94 226
<< nsubdiff >>
rect 36 609 94 646
rect 36 575 48 609
rect 82 575 94 609
rect 36 538 94 575
<< psubdiffcont >>
rect 48 226 82 260
<< nsubdiffcont >>
rect 48 575 82 609
<< poly >>
rect 206 634 236 660
rect 206 460 236 550
rect 145 444 236 460
rect 145 410 161 444
rect 195 410 236 444
rect 145 394 236 410
rect 206 285 236 394
rect 206 175 236 201
<< polycont >>
rect 161 410 195 444
<< locali >>
rect 36 609 194 638
rect 36 575 48 609
rect 82 575 160 609
rect 36 546 194 575
rect 248 609 282 638
rect 248 444 282 575
rect 145 410 161 444
rect 195 410 211 444
rect 48 260 194 289
rect 82 226 160 260
rect 48 197 194 226
rect 248 260 282 410
rect 248 197 282 226
<< viali >>
rect 160 575 194 609
rect 248 575 282 609
rect 161 410 195 444
rect 248 410 282 444
rect 160 226 194 260
rect 248 226 282 260
<< metal1 >>
rect 0 662 330 696
rect 160 634 194 662
rect 154 609 200 634
rect 154 575 160 609
rect 194 575 200 609
rect 154 550 200 575
rect 242 609 288 634
rect 242 575 248 609
rect 282 575 288 609
rect 242 550 288 575
rect 149 444 207 450
rect 0 410 161 444
rect 195 410 207 444
rect 149 404 207 410
rect 236 444 294 450
rect 236 410 248 444
rect 282 410 330 444
rect 236 404 294 410
rect 154 260 200 285
rect 154 226 160 260
rect 194 226 200 260
rect 154 201 200 226
rect 242 260 288 285
rect 242 226 248 260
rect 282 226 288 260
rect 242 201 288 226
rect 160 172 194 201
rect 0 138 330 172
<< labels >>
flabel metal1 s 296 410 330 444 0 FreeSans 44 0 0 0 B
port 1 nsew
flabel metal1 s 0 662 34 696 0 FreeSans 44 0 0 0 VDD
port 2 nsew
flabel metal1 s 0 410 34 444 0 FreeSans 44 0 0 0 A
port 3 nsew
flabel metal1 s 0 138 34 172 0 FreeSans 44 0 0 0 VSS
port 4 nsew
<< end >>
