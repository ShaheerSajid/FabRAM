magic
tech sky130A
magscale 1 2
timestamp 1702392439
<< nwell >>
rect 0 488 394 696
<< nmos >>
rect 94 201 124 285
rect 182 201 212 285
rect 270 201 300 285
<< pmos >>
rect 94 550 124 634
rect 182 550 212 634
rect 270 550 300 634
<< ndiff >>
rect 36 273 94 285
rect 36 213 48 273
rect 82 213 94 273
rect 36 201 94 213
rect 124 273 182 285
rect 124 213 136 273
rect 170 213 182 273
rect 124 201 182 213
rect 212 273 270 285
rect 212 213 224 273
rect 258 213 270 273
rect 212 201 270 213
rect 300 273 358 285
rect 300 213 312 273
rect 346 213 358 273
rect 300 201 358 213
<< pdiff >>
rect 36 622 94 634
rect 36 562 48 622
rect 82 562 94 622
rect 36 550 94 562
rect 124 622 182 634
rect 124 562 136 622
rect 170 562 182 622
rect 124 550 182 562
rect 212 622 270 634
rect 212 562 224 622
rect 258 562 270 622
rect 212 550 270 562
rect 300 622 358 634
rect 300 562 312 622
rect 346 562 358 622
rect 300 550 358 562
<< ndiffc >>
rect 48 213 82 273
rect 136 213 170 273
rect 224 213 258 273
rect 312 213 346 273
<< pdiffc >>
rect 48 562 82 622
rect 136 562 170 622
rect 224 562 258 622
rect 312 562 346 622
<< poly >>
rect 94 634 124 660
rect 182 634 212 660
rect 270 634 300 660
rect 94 519 124 550
rect 44 503 124 519
rect 44 469 60 503
rect 94 469 124 503
rect 44 453 124 469
rect 94 285 124 453
rect 182 448 212 550
rect 170 432 224 448
rect 170 398 180 432
rect 214 398 224 432
rect 170 382 224 398
rect 182 285 212 382
rect 270 373 300 550
rect 270 357 350 373
rect 270 323 300 357
rect 334 323 350 357
rect 270 307 350 323
rect 270 285 300 307
rect 94 175 124 201
rect 182 175 212 201
rect 270 175 300 201
<< polycont >>
rect 60 469 94 503
rect 180 398 214 432
rect 300 323 334 357
<< locali >>
rect 48 622 82 638
rect 48 546 82 562
rect 136 622 170 638
rect 136 546 170 562
rect 224 622 258 638
rect 224 546 258 562
rect 312 622 346 638
rect 312 546 346 562
rect 44 469 60 503
rect 94 469 110 503
rect 164 398 180 432
rect 214 398 230 432
rect 164 323 180 357
rect 214 323 300 357
rect 334 323 350 357
rect 48 273 82 289
rect 48 197 82 213
rect 136 273 170 289
rect 136 197 170 213
rect 224 273 258 289
rect 224 197 258 213
rect 312 273 346 289
rect 312 197 346 213
<< viali >>
rect 48 562 82 622
rect 136 562 170 622
rect 224 562 258 622
rect 312 562 346 622
rect 60 469 94 503
rect 180 398 214 432
rect 180 323 214 357
rect 48 213 82 273
rect 136 213 170 273
rect 224 213 258 273
rect 312 213 346 273
<< metal1 >>
rect 0 662 394 696
rect 48 634 82 662
rect 224 634 258 662
rect 42 622 88 634
rect 42 562 48 622
rect 82 562 88 622
rect 42 550 88 562
rect 130 622 176 634
rect 130 562 136 622
rect 170 562 176 622
rect 130 550 176 562
rect 218 622 264 634
rect 218 562 224 622
rect 258 562 264 622
rect 218 550 264 562
rect 306 622 352 634
rect 306 562 312 622
rect 346 562 352 622
rect 306 550 352 562
rect 136 522 170 550
rect 312 522 346 550
rect 48 503 106 509
rect 0 469 60 503
rect 94 469 106 503
rect 136 488 346 522
rect 48 463 106 469
rect 312 444 346 488
rect 168 432 226 438
rect 0 398 180 432
rect 214 398 226 432
rect 168 392 226 398
rect 312 410 394 444
rect 168 357 226 363
rect 0 323 180 357
rect 214 323 226 357
rect 168 317 226 323
rect 312 285 346 410
rect 42 273 88 285
rect 42 213 48 273
rect 82 213 88 273
rect 42 201 88 213
rect 130 273 176 285
rect 130 213 136 273
rect 170 213 176 273
rect 130 201 176 213
rect 218 273 264 285
rect 218 213 224 273
rect 258 213 264 273
rect 218 201 264 213
rect 306 273 352 285
rect 306 213 312 273
rect 346 213 352 273
rect 306 201 352 213
rect 48 172 82 201
rect 0 138 394 172
<< labels >>
rlabel metal1 0 662 34 696 0 VDD
rlabel metal1 0 469 34 503 0 A
rlabel metal1 0 398 34 432 0 B
rlabel metal1 0 323 34 357 0 C
rlabel metal1 0 138 34 172 0 VSS
rlabel metal1 360 410 394 444 0 Y
<< end >>
