magic
tech sky130A
magscale 1 2
timestamp 1703656013
<< metal1 >>
rect 985 806 995 828
rect 831 772 995 806
rect 1051 772 1061 828
rect 1079 110 1089 132
rect 831 76 1089 110
rect 1145 76 1155 132
rect 2179 35 2213 1165
rect 2179 0 2301 35
<< via1 >>
rect 995 772 1051 828
rect 1089 76 1145 132
<< metal2 >>
rect 0 1057 53 1165
rect 995 1035 1051 1045
rect 995 828 1051 979
rect 995 762 1051 772
rect 1089 909 1145 919
rect 1089 132 1145 853
rect 1089 42 1145 76
<< via2 >>
rect 995 979 1051 1035
rect 1089 853 1145 909
<< metal3 >>
rect 985 1035 2289 1040
rect 985 979 995 1035
rect 1051 979 2289 1035
rect 985 974 2289 979
rect 1079 909 2289 914
rect 1079 853 1089 909
rect 1145 853 2289 909
rect 1079 848 2289 853
<< labels >>
rlabel metal1 831 772 865 806 0 SEL0
rlabel metal1 831 76 865 110 0 SEL1
<< end >>
